PK   �eX	r+�  �Q     cirkitFile.json՜�o�8������2DIQyܽ=���E�!Z�a�+�M{A��#��?b��e�]\���9�!%~83��>F��l��h;��ݦn���Ytg�����̢u��}����.�z�������E{�n���ȴ��X-�2��X/K��Jd%+0�$��	�UZ%Ϫ��Ţ���y��4-�s])�Y����5�t�ꙣ.:�t���H��Ԯk���䀓�<��%N�p�'�8y6B��5�v,8M\䘮���!WC.�\/I<C"ϐ�3�AP��Xr���a�cS�z���#��H�9�z���#C=ϐ9� �l������?@�H�`��i�;)�U�!w'�O�{Y��hD?UU�Exự0)�x/�L0a/SKy?����I� �A�%!�"I�(/)�M�%���&W��^H�+t�kb4��ѬF���aF�0�4�3��S&��!�(��P�i(�4s�9Ŝ�bN�yF��i(��� ��h(���b���)>�����[�7v�wf����^8���er���r�&��x/���E^&��x/��KJ�E�x�hإ�$F��"`D�f0��aF1����P̉"9Ŝ�bNC1����P�i(�4s���b���
���b��h(��bW�7�K�;����Kt�g�C��M�^����]i���&�Q�V
l	Y�d���g˥��biR�D	�|r|{��?G�| �yڰ�X�S�f���j��\�����\O�B�Kl�M.���>qg|{���;{�~v+�4eh�߸A:c��_��~H F@���޼ۗY�o�~HL�s��o߇���/&G�K��Y��`�m@�d�!X���㓏��m��O���۪����ۺ�F'�~��ү�q���+w#pM>�~�!�s�Q5FH�@��^"�
�O�z��g���3�i�e�a4��p�%�agXFR��t8b��zlQ��c�G�a,��)�rʱ�r,��)ǆ����O�$�D@�XK"`I,��%v$>͢��.}��<n|�=�������c�O���6S��h���H�_�~S����~�3�3��fޜy��@�yk�͙��Wp�����^���{�
��+�W�W�W�0$� � � � �p��-~��U�����w_�?�����Ǩ����d��D=1�;l=�q�6��z�Q��,��3uS�����{;�١��7��&~��M�C�Y��egM�l��;����W���7� � ul�B���elD�ĦТ0)�%/r���?��͕�.��|�v}�*���	+�LAƙR2�2KR)��9҂tZ�n�Ft{�6�4�q�=o]w��v}m}���ek7u?<f#���Dkƞ�,�'L���G9�~ߕ��T�U&K���n��xiM,�V�,�ݮc?��/��Y��go�b�hR,�EmW;/f7�h�wE�+�|�7R�ipc>����K�c-ɘ&գq���tԛ�B6ώ-\���CK����lL��Q�ՈQ�jب&�H=����!yz�DpJBfBBf\Bfvf!�BfvBf�Bf�Bf�Bf�f!�BfCf,CfFCf`CfzCf�f!�CfȅJ���� ��C���?�۲n�a6bs�s���?�_7�/̝���������}�,�lV[��ï���e"_Sl��%���ks�>�o~q���ʬ6�5nl����˕ݿ�ٿ�ug]��]�r��4�����ݷ�plv4�����׶!ʫ엦.Ձb w�f"w��8N~̀IR��m&ӸdEkS���I30`�&?�*�M�ALH~B�@)��@���Z^��|G�~�"'P�C	I&��Dd^��x�'��R��܋K����6�@[ߺ�q�����V�� s-a؆<�e���Z��"������;o(���R���W¯'��n�w��y_]w��~��ÿ����b{\D�7z�����E4[8M�_�ͻrhz��dpf��&nU_�y�@96��W��ۺ�M78{\,�/F�W׾�ð�7�ݫ���>���$�y�Y��$���-����V8�x��V�O���Aw
��A=J�� M����I��J�L�+�02���++�����0@��)bt Q F�����I��?�V��\%�S>�j�Z_���*���sJ|8a�I����'y@�Z�(���Q�N�d�t}���Y�lJ�9���˳z�z_�fz�ծ@vE�cj3���c��\nV?���z{�Y��I��_PK    eXǐ]zd� K� /   images/2a01d32d-a809-4abe-b296-5e1ff191d201.png<zUT\���n����6xp'�C� �� 	'��4hpw�����ǽ���sN��N����]�j�WW���I�	  p�e4  �������u��Bp��$���< h
2��^&'�h�����*kE�g3"��n2'�5�k���}��z��k��Qr*��zQ�E���P�AU.%}�����	�;ޓ�k�EA�������5��Y����� w�+H�UhQ`�����	�dC��_'$�Hn���o�)B�х���Զ!b�`�[�������߰5��:�r�v��khL �t/�����v��K_-)��i7�8yol&�ө�������;�FF;����d�^#��D�a��|�����i�2���O,i�B�K)����SJ���	�d�`�-ǺU.��I���_�a+^��G�+�X�Ǹ��K/R>2��W8G��R�%�.��*ou�G��/�H�9u��{<i��'�G���'�*KR���k��n3V �6\�;l̊�n��K��x9���r���9�/�J�h�~В,y�t��J����L��H"ˊ��r�k\�}ff�ƟgVH�a�
�q�,T�l_V]z��)���<�#=�B�6f�z!�]&�5��.;ޤ��V�������r�{�n���������)Y�km��~��$�� �gz�����̸YN�#�f��x��~z:ٞs�t4hӨC|rS�ǅ�9?�UFr��?M�?����|�>\�5En�$GF]��O�=�_-;���>|֧=�!�����X�38x߹�s����SǮlћ���ۂW"K��� �r)��pﺐ�9��_��vw���ֶ�NW�Η��G�ZVe��?����Qۅu��|E�켙Qz����̮�+N{�%��U�ݪ͚D��L���Z"k��Ǆ�J��%�k���< �z1�*���Jy��DͶ|Z��1��3��
�ٴ�d7��[�7�s��y�j�sL�kH�\�o���H8��t:�5<�+#��6?̮>`�H��&)ο�P111�WwN��ڧ���*$0&}h���:%��d��d��۱�5���a쳨*����'�A!�+��G3�)�t��]E�0G�4|�@�����]�=�'n
3ާ�����0c�oi�-3g_����Y��8;q�t������Bt1pVc9#⣙�tӷu��p&��������(w6>�T��i�
��i�|4��@k�lHش?m�J���敒9DX�\N�(�
<B��T0�+k�.e���3��	��!���*���l������Fυ���w�o�Yz�]O���)3��P� �������Y�E��a�k���VUq��in(��L1q=�5��s��,'{1��L~ ��d���<m�t��n#���y5��ξȸe�N<�B�x�h���0M�}��]�C����4�|�ʯ�;~�\���<"1F��0���(����cCgK���;cqC�d�����5IZ�ln���_�Q�����Wnr����Y"�ٞ=�%���������g�)~-�����O���%ȈA�����cRdR�}t � bn�����8U����d��>��i�����IN�_?!�}Â)�ӃfN�j��z��{	�E/�vj�-��gBrh���F��FX��AꜾ��h���G��I[�l�Dds��if+�Ṳ�q��>�l^kE/ݧe��>��߀e����·\\�������<�!���GPeG']4��k����F����?TE-ݐ<8'k+s�0��Ш�����x]j��U`C����]�D������/��M�'��⚊�y��26\U���~@
ش�+K�S��CZ[w��`n\���p�A�u��h�x��fcƷ��_�c��N��!/���*~G���Le�Aċ��
2����!"�0m�Oq�ّ��o�v��'���=�r�1Fحt�i��BC���يO��]sB����n��@����1��VМ��K(�}������	�}�(��V���%t�p��UI'�^�P�7-��K}�:>bk������Z�S�W��T��sW9}���}#�>�~�����Q�bР���bBt�rF��Z%~2�c�����������B�!
ؙ��μ��pu�S��Ɏ�PF��Yۅ=�5�[�e�J�$����sC�(�"�tc��2'v����%�A$d�9�z�����w�TmE��꽍#�)LP-��>#��W�.vw6=D���
	~ �l��"�n=w����p���Q��Q,��j��LK�7�vU�6ϔKX����{�����3fݥ�VH�����W�+�s�ȵ_G���fz�+L7�e�8�n.�Ґ5�2���#Λ�N&-�Y�P8�CC�g��|-:_,��{���4�zb�Ð���Qң��P���I xP��� �@��pR�=�� �Pm�3��|��l�Qd��5чV���A0�}�v�{wS�� ��jX �)�s�e��"E�"�����kF��/Oi{ �n�*$�<氿>�O��4Hg_!1�fc�U�8�c��ke�R�9)y�(�6N��T0�tUi�ܜv��]�e5씪�ٓ�f��%��,�b���Ǝ��/CJ����zd�(���!=����*$�G�kq߄;����s�r� �QZ�V��]��zE-s9��8���ɛi��侮��չ'~�A�s3�TU�����#�(�G)�-�K�=�m	�S��S5u����U�ܮ��T�}[n{���H-�Yc���~�ը��{�����=����\�����3B-����RNB��_i�J���8v;*k��g�ܶ[����AU;F�$]���2��.dA`�� s�w��8h���~��x�~?Z@�뚸��\.�pD��O�����h`���@��X�~J��K����|O�_�᩻&i�1d��>[�7�:�1�6]�bW�RC�E|6"4|���l�tn�#]��u��J���o������a5��/����o�{���-i�{nu]W�; �z<	���_��(�֫���F��nM��d0��۵�@ ����ˁ�2�v�t�Oܦ|k)>��+4� ��=��o�/�%��~���[�92��/]/{N�ק��}���ވ�&���jwP
��dm(�AN���z8����%�Q�Aܕ�����@�/�U�s��D���gK��N�����WL�G��un���!���O�U��f6�2�*�?`�
ui����^�q�*_���ٷ� n1M�	O�����Y�|^[��~�R���_1�~��~��|�;��bP���"�g��訬��b3,{tt��� �O^)1aw���rнvZ�q� Jʗ�)�5�+0�n��y�4$�5���Ga`�Y���H
e�5F����~<��Z����s[�a?����̴�P�^{���>�r4�]��f�+�l��1�tߖ��o�W�{q�����0�Eد�?�$E����.��;w5�R,8'T	�?qepF��zf�!�UX.�i]Ͷ��S�/N��{i�����Ǎ�����sEc�7Za	����B�	O͐�Ւ����=<J����fE���s*�U���2�
�'�N0���ߝ���m���A��՝~���~���ߢ~M��ņi��j��LŊ�k��x���f��{�s|s��Κ&�K�-z�$/�g~���T�5~*�+�gr	����>a�܉b�*��M�J=�Ӊ~��^�7)z�f_��$�����5������o)�Fp�MQ��N�B���u/<��ڬ:z���='��?���J&�:��8����U%���� Oc1c]�O�z�h�/��LŶ7�h�\!�~�7)�II����"�����S����y�J�M�`���]�m�MN{�xh���Z�s��ƚ�u�������/�D�r��s�2�`S�s�7c�>�	ճ�'�}S����Ӥ$�����J���WLV�����5��t�����K���x����q�kd8U��4�?��?�O��¦�T��_�L�:�,W�^��l��H`T�3��P7d���3�����(��"����N(^��S�Q���+�K��������⼋�Ѓ%��	�y�9����݉���~�}oܴ�&k�;\$rw�J�`S�����A�ۯ'�u��n�|^ú巏�㧳n�k`�'��S6fV�x�M��� �����v0�ړ���*"�9��
ٸ_��`n���9x~ �e������\o��:���7�%&^���k�?�,܉V/�B~���Ia�3�q�=N ��t���=������-�dU�w�$c%���>~���O����c�)�#�O��4���w^�H�R��I�Jq7�@a�E*o��u"�E�F�L����̬m���M~���;��J���S0HiJ�2���lB���b�����OW�Lfz�g��T�m��ԏ��	������-����;��Ґ�(H�I`�.[�%���(�<Pr��8F�"01��>�/T�PCS�:�b���(x��[?��I�������_��5O�)����� �=�m7��H�y���c!#�Xm�p�P7<`��EPD�����Cm�?!���[1�.��^���l����p�6� px:v�ⱡ'8T�,���r	��X?b�@��@��&:�̛�L�*�׹��4�J�e$=�{�
:~|g����|�!������:N��$a+�9������*Z����j[
Kg�����}Eze�j�lM������B�Ϝ*�I�@=��6�/�N���D�W5m�}0�� {a���W�q=?eHP`9�!�����VQ�?����*rJ9�q`O,��L�H�����������K�ݱER�a��@r�ȴy��P^H��`P_��u�������I�U��bD@?.��^�Mv�wN��n�p���[��a,� ���B]X5���?�qzP����I���m�wcK�lE��5���OYh�,e:+���靏b�HA�^eo���ybW5X�9��YBޑ��T�Sb��{ni��z�p_
R�o�4pc����i�Z,����`v�d
ėbv�W�!�4�wj�N�*���y���3�A���[�/��&���fX�d�oC4�
���+2Z�B��$R���
 YSu��P��G��L�m�*�+���mVp�]V�ix��%`�/�]E�-"�w��M��< V�7�ȣYL��k0�P�g#��ڌ������`~o4�c�0q#Y.�4z�������e��� $4����㪙��f��zǕF�S6E�)�+T"?�Sq�P�ߚ�(��l�j�����{��w_W  ����K�ru���-!fjm��18��="K����ڿ���Q������k�uFDgD���?j�KmTk$J��	α �X�����$5�1,7��~�����d��]k�����)p�\�n��.������F�{�jƎF�d̴���mX�dvg8�����3WHC__!�ԫ�[��[�	B+>E�2��@��3h��5���'��f�}J���zF���6>/M�9�ϝ��^M��b����[�j9��9-��*����Uʥ�+M�J�m�l�U���&��7�䢺����P�b&�.��_�1�N�y�>\�z�9.[	���ǫ�K�<�����Im��:�m��?�+#'?Q���ǟ� �J��OXgv�>���{9��=/q%l��C�f�:n9�*)&]��'�j�LNz!Xkd�&me�<Ԉa�J���O'��O@��4h�wL���ZYխ��xQ�C3�.#QT��R���ٚ\3	\Ԥ���ے(�����_�h�
��}c���U��]�_���Zj~�jr2eec+��d�B�:B���I��^�$I�#� �N��0�fe�q��gOT�U6���� �f��]ۑ���}\���b����:o��ɗ���fb���\�茆�ژ!��Y�x�������P��?8����nch�i"���շP�Άh�'eP{��̻����{8i�wa^�b�qw�vt gls~n�����@�7�JƸգH�_!�����t3�V��Ȏ��T���|������� $ ��r!�8����Y�X��;�7�2W"*���+]�Ի���2������o�P%����C���ҍO���6v��V�)�	����X�$��w�<�l�/�}��h2ǟ����ӛ}�K���	��Ҷ���]�(Wgf������Ѓ�	�zmmu�%T(����F�sY1n�O�+hb$�$Yon�w\2��Y0��r�9������=m��������h$���Ğ+}���ǭk�z�Y��Y�+Ĺ&5P:���H`�%r�|��%�sݛ�t�gw�i㊗��]S�t�B�A�g^M@�'��@T^$�_�l� �x8=�"=M���w�%Z�2�Y/��O۩�'u�:V�2�U8֊���c�v��C[Y���:����0�����Xшo_�������Q��<���Lhܦ$ad�{&���w��E�<��*�!H�u�|�^��M%AH��7gk�8��%{�� �o�̸�)�����	��O�	���	����)���@�����A��A��kD��>�t�m �D��8�A*�m&e�J���<��c��U�I�p'<��]�+�Y.ܤp+����MB��~���=�cN�3�������m\�lkB����W]�ǩ�P`ӼC�gЈVֽ�&���b��p��.�<ߟa�/ۣ�6a� q�L�o�A�L�^t��y~��e���������?B���:��?#;
_NS4{��/)N׫��Sl�f�'M�2�X����<!���ݻ�{�F�W���n�'6՟�����6�̤N��t1h����e�j���^�d�"r`xC=By��K��L|?s�����卟�h�xPuR��r�}��nc�0;Y�m�	!8�A����&���O�ߜ�)x��!2�:������=���7{P-h����bШ�h@41+��	`���}4WF�I��k�!WhS�L���}�9��"v�[��m���Q�6IU�m�gY\CT���ǥ�ĬG�)B�Gs-�D%���єj7������/>a��/�:��uA��
��Y�3`%��Rc_�x�3{��d�Щ�r��p�i�XV,�L�ڨ.�[�n�r0TS���$�'�x�����]�	O��w�\v!�FFDx�^�͂l���|X&N��3���P��^|��؅��:ϑ�\ ������ �Yq���-����q��C�J�z�@�7�+&mk<�e0��~��t!�b.�OY����R�[̘z��p�&}RUm/��ҿh���ߟ��/I��_p3$��#��Z��&'p���ɴz��o�s"�X2�)q��z"O�)�.GP��X)m_+����'G�u*Tŝ�kHҭ��.�mȶ�nX
�gg�P|���,�%:i�.�"����i ���3��qS�W����4�R� �v���esCd�~��w�.��u"�=s��bv�NC�  �s�0e��h��˙g�h�� ���8x*���Ծ	���R׊�5��᭦�{1g�jֿ����_�{�Ǥ'lRc�z�#0-���Q�4�41~��-���)��.��������jFZ}RJuq�L�*`G����Ҫ�Վ���r�J���9�ի�h�������m)b�/u��.�<��6��2�BM��-������s�O���U���~��͙/�dyd-����[�Kq�mXM{Z�/�] 52�"�T��-f�\����J�k�V�k���U ��C88/u�H�Ġ�@��y��n�/��(�Hq�"���ȗY��ea1B�4lOeu�g�kJ����s��͡�8��"�5D�{�����+05�L>M@��Dy�e�l�I
�ȶzw�����A�����a��{o	�=@U'���Sd�^�����ytz_�_����u>̷Iw��mћ��܅
�l9O�sF�����|5�:���	{V豝�A9Z]Pg�{��~�C�Ƴ*������1����3!��(>��S<WcQ+q��c�վ.Cy�qP4.�x��ǈeh^qU��w��Ƀ�a�rN�d\�%�3�D��]��	� �4��fv��E�c��6�^1E��v�	��_�
�@���r��l~��h��{�Ag RP�~'�r��p���1*�W-�/
�(<Ȅ�ʐ~�Bu�켓� ��hx'S��A��6;F�q6�E��>տ�fUZd?z� ���H�E�9,�GE��S��$]/�Wd]z�{��¹��Ju�1�|�9>���U#��E�����?��R!v��%�
ٜ
�hE�"n�漱����5T�-�ٖم�ݮ,)J�ܨ:n��$�A����h������vK��z�GS��+&�J)������z�H�T-�Dج�4��3�LN9�u��`�y�
�>^P<�I&7��/��%:��F#���oɒ#N氎��d�۹Zs>o&�4�#�'A���)�f�*���#<�Ͷ�m�w����?d[���8��ƻ�U�ET��L6�J�D�:go����&��[����(�� �D�E����7�y�P��;�Ks��kn�m�*��r[Q�Q�"dH� ՙ��t�_2*(�:��z�n���B�Qi�N-�;B}�ژ� l0ZVnD)���
ǐ�2����[�;[�E�E�,D�Õr��,�%ܸUx%��&�H��:�e굉������'#�X<�7B2�����R����K�Xoo��&,�T�1(s�<�hM������+W!R�g.:�O���";#o�~ˎ���a<\�{�iP��ś��<3;�:�=��nzg8l�aC8%Z�*�ŠÂ���o�����4�&�·��X�*�㢶B����츉�˧��lo�a:�3 ����T�;�)w��C������R������y���Wg����.�n�&<�u�^���rr���zȕk�8�|S���/�� <�w�L�Y�;ӛZL�)D���k�V�����\������]�I��ӹ0a�t(��\�j!̾��\�x�?�G�i1d�T+(K�<I�,�i��w}���k&G&���P%�D�Z	��5˘�����g4c�<�۔c�;0)S&�K�;�����<���Q��ϻ��ZTt�]j��J���l�}|��\��UC�y�Z[�Kժ!�E�Xhucw4%\2#"Al|��ƀժ�.{���q�L�/E.TC�oI�Z�x�b:UQ�1�!�)�5����DšR�*��_�z��$[�)���M��1n������cbP��4��
h�����V��"ǜ�?}Ǜ���߷ߨb���Ԇ)#���j/�����ٹ.��>�����t����Ƌ���M��V$k։�$[8�#�7YYX�z��q�n��L��Ɵ��.�?��>B���s�8l\ϧX���ZBb�$�]�8T�nLm��'|~?�ʝ�K�����-��������u[�X�6�Y����[��K�m�$)��Ȧ[�'��c��cɬ8f�7A�W^�|��p����?"�WՈ[I�$�2�w3s��a.Xl�u���CPl鍍�[���͂Lf�����Px�Z�������;�4<q(m�o����+��%�w����:T��=�9J�4�[v���@M���Z�<+��#	�Y�\gzj���;��%W�7���v���Z�����gaG
&��o������uo��\�*�Ci�Sd�齅�X�K�x]~�k[Ä�������pa8��'���;����J]`�}pF�$k�aӿ�]�b&j��ZHJ����[�Nj[��{u{����m�s���N�Y��&ݙ��qw���x�2�Ѭ)��W���g1`KzI�-nzX���_N���-�#�?7j`��r�/[�D���\>�u��L�Z�13�o�B�9.���h�4�$i2Y���"�����,C�؉Υ�-"� ����u��p���ꢁ���g@�������۱�`�=I;���&j"����NmJ��am٢�2WP�&gr��#�2�D<j H�(W���B=]��?���Nf����/N;t�"���t�}�tOF`��S�+jRԸ���d��G�����i�H$= %Z�}u{c	M�0];RJzD�<S���u�v�Q~)gʎ`B$��Hf!��+Ֆ^���̠���_=��8ABL���Bq��zb���R�W�rImK��� �WpK �=��c��I$��3��	�Q��_���z5ʥ�4辉@�:,J��'&bY�A`�xr�s��sm�hD�&�+9�O����tk����q����Wr��`~��� X`������֛KS��������������)��ő�x/eV�C+,v� ���*S��yW��<~ �4� ?�$�i�C���V��w��`�����Ub�`������Y�%��}	H6��P����B,"�G6��xW�C����'x�H�T�����e��W�<7T�GN�����'[�caE~Ks�3�JGN��t9���3M�_Ռ�-�y�;o�S�������zC�c"k�%���6� �b�e��x\#�� �q�|��9�s�]��eM�fV�E�/��ą?&s��:U%0Q	e���F'�ڇ��U';�C:+��wބyMy����*Y��|ǫU{L�e�,�9e&�n��«4h�&�4Rݴ��&�K�N.�%�Z2����\،�z4G����lk/V�E��e�s;�
U�����du�`g�sҾ�$�9	\�������beJ�P;ߣ�aml�P�y[�#��������_�a� ��ƶ�s���� ���n�
��	���nҠYD�OY�aM����y���u���>��f<ݽ	N��Y�&�����eq���{���9O����(���&~M�� �Ѓ!��?����*��!Ѷ#��!Q����V�C,H6�7���0]���ϭh�h�c��9���{N����?�����h� �z:57Bb�Dy�D_%�8HB���Ys���ęS[JsY���@A��O�^&�9�+�k���e��(�n߹De!*���-�a��58��:�C�~��p�fiF�1�1�1Cn�������DJ�m!лTWN'�,����8�>���A�
1����c��񥧧��f2����e��I��������"���=��!�� H���=c����rj��,����|6m۰�8!\˱��Zo$�;G9����mmy�cm�^�QgHTxIƕ���N�8	����˭�Uܐ=�N�>le>�|�i�̀�ާtt�x�7�u�<�o�es���"C5>��h�c1"Vo�l|M*��q��wk`Q /-���$�y�w1�@�����Y+��]w/+�� ,��s�׺5)�}5~T�a��i�o��hH����?�b6;���OL��5�|C�i7X�<��Ϩ��<���+?7�kao�`D�)@Խ�ː��l�?׿��G��_֎�A�PAD��Hj�#-��-�xi��3 �'�H�H�Y�-�"b6�y9@��=��zW�A[O����P{f�)���*¯h����3�B٦_)�4/�E2m	?�M2�h�#d♍�L3�����G�7㏕2P~.�3N	E����������ܝ�B�y����yO�TA��z�/&���BP�d���u�;`v_7]|B�I�]8��Xn�2h�87�{݀�%�]#��;�����ʈ�0bA�� ����#i�a���D}?Gћ*ɻ>q4_j��^q!��?n8x;WR�@!o��(��B�Z��hh���_�|��§r�/Y�(\���i|���S#M��5��O#m�@} 
ܠ���E5�������'x��\���'�y��̅y�Ɠ�ѧ��d�>��*���&�Q��tI�_1���3�`;������B(�:Y�P��`�<[�NŘ#Ή(��op��Ѥ�y��M�M%�j�w�Xۘ7֬`����R,���/Uk��0z��?���wD�0�V�~i>�"���/W�S[�?V�DHBzs!��5�(v����\������fDh�PG �������xۙ�����
�WR�+�j ����x�Tt��p/�$���������ĉ��;	j���j �⎸���ƊweI����	��k�X�13�\��ݓ}�
�_w_�����=���HO��m�v-�S�-�U���8I�N�����Ln�
ɭ�s\d�ɸi��`;`�Y[�Gji��ґ5�*��o�!�C��)�������p��a�z�Jز^%ʔ� �� �.��;�X�I�Q`�G
�y*�xf�3B��C��@���%"�<>ܜ���7��MƮ��b]���o�m₌O�<�A�@�g�Z.�u1z�����D�΍�u�S�fo2-���I^�R��t��0��M����8����H��h�ff�8��<�M���"v��Tؠ���f�����z�՘C��Dٟ�xɡ�oe�����paRD��W��1m�����* �k��<�.� �wo��.+03�W���[���bUQ�g��,����T����џ��l�-�+P�	�x�Ar1ЀBc��1���ˏ�wJ�� p�oN9+:@���8��RKbBN7�N+ӿ�crrO��[�=.�w��d(/fj�lV��&X�;�ϱ��ຉ±��@�;�D3Y�bCY�L�)��@Pa��6*�S��[d=#�["���R74�����&�֦$I��1S�d��[7�;t�]t�^��7B ����q��u�N0,KS�\�X�(�8��C�q14�*!�B�^Ϧ�������ę^I�~\,ߦ�Sǀ |,l���[��!��z��[ɲ��JS2��Ԩ���L�x�����6>	;�cYX�S,od�HK�0�i��ᓎ���o�m�Z/�ӻO-f�U�F�c�7m�����	����;YXj�̓(�$���H17���x�ӻG�.��Y_y�vv�	�tww���mrTRFq�+ι��nY�tj�?Ŗ���uY�{砑y�o��6�1��"��5�7#��1Yʴ�	��ϙL�x��+Q��&+��Z���Y�=�3�֖q�K]�*:I�����$!���t�Z(q�oXI�jdB]t�0 "ÛKΊQ߅��	jɐ�>�!Tz���}b�d)�`3�]��m�Łs\��=��=��e��m슧ў�  ��vM��*�Jҧ���'C�y\F��F�*?r9;�uM��I -v��R?Zy�">�IY�s�ʍR�=�-A�<�?ݓ���)�P��vX����{��1x̤j��Z�c&��O��{�j ��c>�4wp����Db�w]~��"�;j4�^��r7W���t:�0@����;y�o�/�xzX«��J�3b�v?�
��Q�^n���8��8  �y作���5H�TT��\U��XNym�3�����k~��ƏwC��J�H�Ny����|�l᪑)�=����'V������ ��^7cI�ǧ#[e��̜�O���!98p� ���欕�`eF��E�Y��z���b7�(�)���1Ż������ԥ�~4�� ��$21{P�[��_=��V_8�������%����#
����b�����3?��.�Ow@�^���H��t�޶��/L
dW���_��I�:��J�.pG�}��`�eQ~3>�/��A���:Y9��a��5q�Lpr��;&U�a�6*����.����a.C	��u�ջ"$3"0�2F Y(.R�^*��;��+�E�h�|��7϶��]-��\y5Iư,O��2F5���"oڶ����P�/����=Ah>�j%��9��
ճ�����T�����C1�31�w����L!�����
l�ɚ&��s��c����R��D�<RS��:�wc������W}�Z�ꊲ�ȁ��>���T���1_�~�w�Db��޹A�v!<TA�,^<E��BF�>ZX5�k�~Cd�Y$�
wÎs
f��&��@v���v��s�� �:�+�Β��,��yw�5�xr��G�a*+.�pZ:�B��/�?"��Ⱥ�F�ۋI�,���xs(�0_J�v��;W�3w�-Y��\����������Opr�Ao����5�čM+�ѯ׵�P�^�i|�puc��VϪ� gd���������-�9��ɗU��0|Co+�b�o�2Avn��ʱ�H�$p���5�w?Ұ�����+�
%3�B�q\i�>�8�@��ꒈ�q��G�N�sYA��5�(�"�Hy��l��Dc������9�b����>b&fT��Ȧ2�C �(��g�	�
%�$�襒��QU��Sد
���K[�a���p(2�gr1 (��z�=�9�Ш��&�H��D1�������-��(�".�ءF�� ˋ�و��S�W�P��������m��N����<u��Wu�x����H��S8D�܏�q�;f6�4�v��հ�uA��%�4%5H"���= y�1���������*����Eo\���uә����I�F4�"�#b�k���,��g�f6?�;U}�j{-�W�� /	�x�P�nĠ�
��n'�+���\J��OQ���q$"��$�S�J�8ƳD���C�. ~�o��$8F#��/r>󞆫�ſ�A��>E�~K�;���&����Q�ꛡ?hq_�~&s$�V��Y�|Q%u�i�B��hM0ۆ��"/Ɛ�O�'=��Եa�I����J�������e��%�ҀH���EM��,/S�?�D���O'�AO��g�h˔4�A�\����Y�b�:'͎����'Lc~�3^�D���G_�����$�v�OC��-�����?���@]"��J��<��A�����q�Ue)s	p�HbԽ��w>Wćf�/�u`�JA[w�o��u�����4�%�#�4�.�RJg�-\/��g�Q��{�|�gTN��[�)�
�MҫA�9	���c�W�zӎڽq'�E;HG01���-���+p{
6$����Wo�:��MF���fv��f�4»Őh!�s�g�A�p�IL���c-u�N�����)X'k�ȖYQ�N����7������7��B���R0z��	�:�8F�o���ԕ�)��keO��ӱ�MV�S>po�/M�J��mJ	(U�ӎi�V�A P�N_i{ �H!A����s�;ć_t<!��ƥJ�3��_.�$����E��:����s>�S��<��+��)�/Ma��{qX�1���e���ڧ��G���.S�>&j"��~[�´L��onYu�n˺SG�0����jG_����+��#����ی��N��t�9����X����k���g�ĳU�we,�ڥ��tM�ӾV�{;+ks`�h�K	?��[�U"u��#| z>6m�}��z�]������)��ltĉ�O��I+t\ac&_W���4��-U/cO�pܜ��U���J��ݸog#=��s�Bh-�(�TyuyS�@��{����BES�l0�9OBPqO�B?���5Kh�n�3��B��Ry���ѴX	�
/���w�VB��"��SY�e���t�8'�UG�I��W
ζ��H������#v%3*�k}n�coO�j�g�*ptTN��"n,�W4_��;bª80������[�D\�$�:��Q0����S w"i�x������]������X�-um �}Ko�P�b7�~�3QY6U���P�z��R����<�U� �)\/K��w�L[}1A��9JM����y����=3������_,�[�#�w�Lm��H�wEiV�8W^	;�2�ն�GN臚f��a�>��(چ	�������'���r��~��I?++����<K>j���O�B}iW&�ڶo)$�|�4�۩�;Š)dc�!�j}�vs����W�U2�=܋$ooL��4��+TΡ,݇eC���|Į�:k�5�I�?���Q��o�� ��ٯi�������g�u�&��՝���cL4���{ն��.n��Z�P�䉨�$�P��vzK�r�D�%��U�f�=�Ps�~0H�?�ԙY�����Ȝ>��#|nh3u)�'u\ד3lr̽��g�n�Z~k� �mrXWtߤg�0�xH�z�w;�7)�+ pIJ��: �e�ypG��޽OI׫�H�\(�'���Ua�S9L����] ��J�o@��
]'��ꊆ��Ǐ�b-D9��~�)
쯝!�D�XM�o�����`o� �b_K�_��=�������NQ/�ڰ��ķ�T*�WS�0�s� |@���Q��T�kTJ�$Tcq�?�����=����S9�Z]�[Ə�����?q�.�%����?�Dwǎ�裏&#�p�F�(_Ck֖R�����9ulv>?��Dh�J*�ї��VBy��>8k��2�N�|���5sf�|���>ӊ�U�.�� >f�u�LW^y9u�O3N��2�F| �"5�a�z��gì7H55u��2������?�T���/���������C�a��.����A��.a�ʕ�F�U����w�Ü�
t�Q���ߓ���./��t�J���~��ʶ�;s?�0d�զA���=���1*�#�1�
�����i(p����������ߗ�)e��c��~�q*-]Cy>����0��Ր�)�z�L�8�y�B���T�R��ǐ��<p5)�*���i��/����P߾}��4z��_��W<�x���P���V]�VZ�t%�0 w�o}M	D3��`fa��ul�[_���<�\�p�$����@�^�CѰJ#��B��Q��������~���|�̥р�}��%ũ���f�z��<��^�֮[Eu5���ϟO�7m���uDF-/�D�FO��/���n]����x�*����Abp|>8v�}�������$(���|p�Y����}��E�6��үi�UL[yL/��w�U�6��y�Q$lq�#p��}z�,Rn����䂿��Rԃ/�U�v��m�/嬟�d-� 6e%b��E�ԱS<�
��x+u�`�r��d�9_�IlH���?�<��xz	�q�i�����oyQ@>T��.@\ȁ	��W]u;s�>7��i�TX؅/YĻ$�#%+��d�jJZ^ڶ��:u)�+����� m޴�����iM��j��ch�"|��5k֌��%%	�*/���ϙ	����M�\{���*]J��EG~F�֮-�Ꚑ]l9@U�:*[W�Lⴶ���4�P�+;Ā���9�1 ��G ���'��'�� �����6��;Z��m��+)T���nZK�C����p�x�h��-4w�����A�!CQ�>�U������j���z���?����W��Fz�����30(���ѣa�E�xS80�z|A2<�o��CǮ�.�3y��(�08�4=L��,�mٲ�����8�^�o�2oPC���1�%�/�0��0 ��\D��y�ƏF�:���ҕ|m���(&-_��j됴.E��A���N��������իv�m]�w N��JQ����W��9�|n޴�^{�E:��)�>Y�a-{ư!(�e�__���	�-���#���C�zı���]���.��
P���JgMǃ���Ac�r�F�֮YF��WR,VE>R�&ȃt��o�<o���~D�5	��۱�0�#0aT4���j�.��K=�#����?�����G���V��+nG��䥗�kdz�s�"�t�T[g�דφU[Q��8�$�[n���)�{��٠[YY�.\��Q�F��(���о�m]t�>˖|I��7?[�N�hU�reo���D�)Z���o;ڴ1D	�K7�p+���y�>���|��t�L?�}l�#p�WΙ9�QW�Ϡ}�G�z�^}�?�����)�{��tđ�r����5�LD�A�QUU-���@���ʫh�I� h�>�(h�6<�r�<��s,y�a��T�38��sU,AL��+3n A^���i$��IR<
�~,~���h���޼�i{e�?����O�K��u�_�=�Ye.@q�Yԛ�C���#x�k��o��ϋ��a;�@:��Q�1��ø��&�
GԾ}7�2�H�D=���6�����2k�!ھ}���;��4v�g�}�����w� u�������|����u�d]s�5�[زq=�{�%<�7u+�H�W,���6;�;*�%h�7�(�C�_������^�3N��y�OӺ5k�8�����r��!�Z?�Pv.��%]L�J����?��:��R�n;U�l�bҜ���i�hݺ
*��Fյ�}ޅ����{���w����d�>x�W^y��}��!0����@rA��u����LI�C��6�	~�@�$D�'�Q�C�(C�> ���K��oSUu��� !=:\���7�J$��������i�?�۴v��'N؟ƌ:H��'b�1�<�����d�Cy��dz�9:���q��H��g猷�z+��C�5ft������4�#���nc��*�B���4�d"BK����D-�UUo�H���>�c	2� ���Bk�ld�m�Y���I��'�y��ѳ�=G���6� ��Fh�$ZG��O��舩G�9g�I5U���I2'�u�z�Ek(/_��HY^
��Q����P^�*9�l�!�4�����p}��]v�et�����T^^��@;�� " ��. �C܋#�2�[층C��WD
zUvB����:� =OЖ���ʸ�����S�~�bfgVt�_�>�Y�q��i��8��<�ݾ��:w�gy�5T1o@����H$T1x�l�k�Oe��y�*� �:�;�<*�ѝz�!��1���#/8}`�=��C.L��O<��:�(���5�T^V��!�����C��C�E/-Y���7�8�|ew�i���胏?�pK��>�x�6��7��ɼQ<�d�w��t�Yg�AÆP,RK�U[��r��8"Q+�d�^Г0�F��H�G�������/���x 9^��	��#!�����R��X���D����M�雯>���j
�}*7�O���─px|D^?8��L���c��/W�w�t_��8`��7�?%���[����U�D�Y!Ês�GdL�rN/x���ٷ� α��T��OU�CN}�ʉ9��g_PM5损~��0�í;|�P'��|0���do���v��`��F�j�����G��W�i�F�rĀM6�~��!�P��9�D����#�������z�x���4���l�>`�lauG�M�<�N;�T�ٳ;��VQ2���3G������CAC8�î۷��	�@�g�[(��u xб#�� T]�u��JE/|�����2�2В�g���i���H�8}-��y��L��iS����T����={��h���>�d�@8)�'ڎ�$H�I�'6��Y�(��2qm��R�Cg$�|�53i�hX�6�PR{�N���R�G���<<�˚�W�ʕ��r]�̰XK��
l�f<�D�Ka�+m�}%�0�2&^)�g��� ��&��NU��ţ!WOD� n��#*�ߏ$��j:��{��, &g�M ��eRׂB:��cXY�=��Gh^)hc�n������!�O;�:u*u�܁�-�џ��L��s���^�U�V����`�׏��Z�1���i᢯�w��[���1��T �G��:��?�A,���S�$vk����*C�eu��WL�,��փ����C��q��m�����x[��o� F�!���oLd�|����|�s޹��c�q�8 �A0 J&����^ �-^�m߾�>s��d\mg�yLQ���@ｿ��a$*A�i���z��co����D{x�n���[��7��&/��A[�L}�	���:�Sg� Ε8e�Ef�.y�)�+I�dao0�C�����p�ް�����"�8O���[{ђ�幄�D�ޭ �,��G�^Y�2�������	��l#3J�F����R; ���<d�a�MR^~'�<�p�/Š(�|\���\1̲8h�w��s�,��j�5���!+�|�|��ǻ�5d�`���0)�>E��	�1�H�_,`�eH�P�����4�7��G��)� �	w�ѣG�ĉӞ8�M�3�H�~�U�Ѕ�ϋ��%D"|=p}��G��(�+��������.��w���3�������z&h��iC�J%��1�DurMP?y�v�F�;�S��Kp��xRe�D\��bٚ�����Y`c����r_�/�#�s�^��8�3W|'Z����8�8Ydd!�׽+�,���@�%ͷ$��;��v�eW�FԂ'�+�"���) �c��[v���󥾄 ��&� iJ�E@[ȿԻ@_�x����kQ�I�O�w�}��_J>3E�D2�>#)�� %y����Qu�h;�б�<� ��GT��~��ڸ��~w�oc+�?��G��]��c��ǜ9s�D��_"��%0����!�"E�eG�>GL�E�@�{,ؒ.�	��
������vR"w�ഖ�6����$��a0 �m�F� gܸ���v���D͐ÿ�b��z+}�����/2^���g��#G�y�����Z��cၫ'4�>"�ҧioJQ�f;��B�(�f?�R���������>��:�*����ۧ��L�j�}t�Z�P�|�  �F.�s�'1r�}��/@+�X��~�i�jc�$x�#�
-����E��sJ2.NyN]C籱�H�~�|J�|�� ��� ���Y}7%�,��]zۤo�|��ޘ빂�|?�To��c���CGR
	�L"V� �RA��ku�\@E�=9
�5}�"N��r���!��&v����O�;�z ����pA�0�y睼c�Dh3�;�v��(�`d�1[�h>X� �ʐ���?\XTpe��i%�������a�hDe~T@Z�dᓉ*�������<0T&����@�2R�"�
�P���q�����s��>���O*߾��"���@����j�"ڼ���*D�f�Fzo�'�d�챐��Ճ���k���K�]c�	}&�4�
`�J&�l�dLu�_^�e�B�H�Ut@����:��6�_�r�����
l��,$2�B�0�E��.� Y�t�^��m���N�Rr�>)D$�+�Q��Y(	}.I���`G����+�0hp�	����G�+���@G�7pu+�G^�H!/��F�n�����;v�	����{��x�ͷ�G�|���#.�����v����(ʉ,��C��O�%d ���� �%��HLͿ�c�\�^�I&\&���ŕ�`�֪��)��,&%2�q����ė��q�G�|��CI�!�i��G�d��8�A2RaZ�v)�Z��k��^Z�v͝�1��*�����5�\ku�d��'ͽ+%� @���g�E ����`ӵ^L^	�G_bl�ѩI�����'=d_
wX�s�w𿠦p}�nF�`<ڀk�}E9�3
 $���e"�c�w�L�_��SG��<�h�����˞���~�/���P�}w����x�V1�Ȅ�X��=���~4��IdQs!Y[�s�X�9p�>���y�F�����@�����[hђ��������@�z!�3(]��t-� n������@d�q�$�t�v?��

��5k��m��9mz��U���f��(���D��\�.����f��Ź�q��`�|�ǵ�L��~�v �>Ĉ�E��^����P���6Њe_S<���@�JK7л�>J�����r�	�plk<��L��"�Z�k�a��h��������ݔ�1������ୁ������v2V� }�<� ��y�E�Ƃ$;H</�{8�%���0�b?��1��)���� &;F�%��*#��L��DD)<��(4rd;O(h3�Aa��]��c��㑘���a�d�v E>�z�J�HE��&��7n�rD���C&<�z�N�(�x�����|ҢD
6b��kp,j���+�p�1��9�}�)]����B�!��E��cA�� :�J�CY�kd�(��nW��1.���"�4�6��5|ݧq��G��k�2x�Q�V_���߲ʋ�&a��	m� �#x?�t��P�����~���?L7�����Q�I(Բn�&zw�'\��4����O��;x��V�G; ~�?�8�O�X���� _{��B�SO=œOvm22Q��Ȯ�>F�$�ɵtZ�Q{�^` Zl��Q�M]�������N���0��er�f'FTD}��w~>����4�u0?�s�[ ��믳���_b��/�g���}�a�~��/~� Bd����K�&��v�(ϔ�=� 8j�6�#����H��b��b�^����P"�����JZ0b�TVM.�J���y~���p+J����g��;{�%R<�.��5�,��GqE����x�]�Г���c�1 S��w��߲����;���`3�ْ��)�.���	��B&���̚� &2���|:_=G�(��|/m�\F>���&����B0ОV�*�y|F�*�컌�?}���&��ښ��<s�L�P�\QO^�LLq)6��	��l��0�Ђ�r����x��y�B mF7,$�uY��#*Z��a�9��LP�"`�äǳ~���gM���y�~�I�&�_D��,���]`����{Pp.�{�M��rr,vx6��xθ&+ v�9�ոq��Ya��������B�+�'��Xu���h��)%�{1���t��jN�fQ2UG�L�'�"�7��OI��ӀA#�������@�s�@6�r?��@�讶>�M<v��s�����D���:N	���j�Yz`ZI�_C�ʋ��>lԁU�vݒ�!��354���y.@9��|�h����w)���D˗~�Y=M�Q���Z���U������k��b1(�8���j�hъ�m}��7�A�`Q���1�-0��Ȑ�K.I�'�Z�,��t(��Ď��������f`��O~����#�0��?b ���3�h x}�_Z!*���\W�S*Z�Î�B�Wp���N`� 9�v�L���n�İ8��x1DPǊh��B9��7�a����]w/��=��=�=�-���P�K�����1���$vK$�h��h"�t�㬷�t��`�R��]8���A���ߟg�tFb7esB�8�9��͝�믲3���z&;  �k�uA0E�[l��ؤ�z�����'m��w�2�]�a�.�������$��t�]u:(� �3�Mhcp	e��j�	Z�b1��[N>�E~o��Q���'��|;���TFY���Ę�4�?s��=�@h��U� S��16���x�@� 8A�������>~�\�VB��K/����cq.���(�@��Y���������_.��_q��)������}�g����TԮh�h@���{���
��BH�,B(����X�d�õ�;Eܐ+�`��n �� �yj�̺�)�@�����Z�\�?���v�x��<i,E�8�c�R�&�׿.gWϣ�:���	�n��~C1�_�{����>����_BpAD��E3�>�3ĉ��XY�Equ��
�~2g��'2��9|�%G�\�	�E��#����%�.=�K��m�����Ȁ6�����	��@�d���b$h��o(T�|��f���]!���\����y�C����O$�5�N %�֚iDO#H�4*�q�k;���KJ� $�;$�B�t�E�@��?!�4=?��#�W>��w��~;����?�1�eq�<�{�w HaW�����ڴi������T���x ��1�(&LH{��>�"�	�h<�	8���L9�98��-�]���s.B.�+D���u`�s�y���E�w4���!�0vM�:�,� ���
�t���	\u���'R4nq�^s����#�3(�?�r��������8�]z]��y���ϐaQ:uW�F4�p�iO�BU�d�}t#��ً6���� ����x��; '~YY~��;�` ��Zj�o�����27    IDAT�(���ƊFԾC7Z_���.+��0"|���߷O۝�u�t�xa ��I18
� @��M��c)�iUF�����uA�����y��ǩg�^�9#�hZ�׿���TPX��x�hh��^�S���c�� ȣ��,V��@����5cG��K ��\�7���6j�Е��5���of�4Y�s�-C�c�wh��E`����i��c��;�B"FmQ��ZN�;~��zVO��f���NЏLJ�$bI�s�.��#�Q )C��<^������b0�/]�2c//ڤ�� �sYGd|:G����~N�aQ��g??��mP�o����P=bm��
t�1�g癑�Y���89'�^U�ro�l����-j�b�0����!�9H��Q�<������˧X"ɉ��O={(͂�����Ř�P
�/솤��h�H�'5@р�����c� ��9@������y�^��c���`���7���� p�\�]Py�߇~�;�@
P�1c�a! �ʽ8��&�馛ҁ� g|�Pa�B�kKIP^Ai�3��#�7d�G���>��)Y$|C6�},hX\�N�+�K���E��}�$^�I�w�﹂��硔!���R��ԑ��d��~��?Ծ]g6�r��]��J��rTSU���s�EC�|�wI:8Ѿ�0"�� �3[�n�'��􀓟�l�d��X(L(�x�`� `�K�-�X�w�q�_�^�8�'&�cnJ�ʕ�i�ܷ�&���~���~;�Y=��mՒϛ��%܏z�(TG��Z/�Ȑ�H�J�ᢿ�cE;�/���>c��!T�ѷX�la=x�Hv�D�\ �C�@Rn�H������q<�����������<�'�P��*<_Q>����Ba1B;�o_\[E�p/����!��RAN�y�� Ա�by�[�v�W_}�89_vI�����F��kz'����sp��D-u��P���k)�qv[D�#�-�z"���ǞH�����s����<~P�w���ڎ�$��9��f��3;�Ocm�!�9�W��u�7I�늑�@��ud�\=ۮ�C��l�d[��~�cF��ɇM��p��l��2�!�xSL	��N��|ݗW�� b��DRɫ�k�Sgٲo��l5�=d%c�1*H�={��\]A�|�5UVE8�F���Ѐ��Ͽ�k����q � ��N:��W=�I4T�%:�b��X4` �5j11ax=�i���L�`��w5vH&���ջ7�
 ��~���.���i��;���ޡEc\Q����y�B������d`�Q]����?��ϋk'vH���(hY���C&���}�;p�0�"�0��XH$L��+�
	@�	H�*�7�<�&����)i�q��.�\V�*e/+�ѣ�҄	�ϓ�?�����~�~k�}ߗtB����� #�ҝaT@@ �E��8��1&�0Bt=���â��d�I��{-�W�V뭻��|���[��Mխ�y[��=�Ou������<���<�͟��T��FƊ6o�b�����X���I2�����=wr"�ց7Y���D,��zW���;�|���^�}_(��yԺ{{�g$Pd(��e�d�+�V�#&)zF<�����k^�j��h��3aae��3�Kֈ��8R鏍��:`���W���F(�`<=�i~29��F��UO�!T�x�N�d�h�\���(|3��Z�r��{�x��6R�K:���z�+(�E���qu���(a��r84�g���\t��y`>_�!��0G6Z�={\�%��G�eB���#�g������B���8�	��^�{�ġ��ݻ����QQ�0i���c��*<'J��SJ
�;4yNA�%��,�Q�<��r���;&B=�p�"dyw| r�J��u���p��5�o �չ��g�^�5�������`==��÷^�͛�{y�L��Ț�綶�V��P�YG�l���W�x��{9���fQ�4{
�~�w��<31/�(>Y��}2���ԟ�w��VB�5�f�:W*�-[�,�xa��T��*���l�����s{)�R���)�q3�f�@,�f������wO��'">���k�m"���m[��*L����X�`�KkU�c�a6/�	�S,�ȨdQ=���D�;^�[�z�N��ju��Y�~��^-Z�����y�sx����6:V�F�bfk׭��+����]ҙM��I�}��#"'\�C?���f2��į����#�F��ɣ�C���@D4��v]�M�0�c����;~��qo�q��C�&@
 ��ً�Z@])E�KX�S�XZ��}Շ�"�uP���(�1��@����n��5{�!͟5��A�4Ԑ�p3���<�G���z���|&a��y۹�^�-�(Y:Y��n��Z��iu�9���q��24Hi�X!����Ü������uA�l,s�k��f�w(a�;�B�e��((���n��;za�cHpO��:���6�4��������mOJ�6��ͥ�^��/���0]3%h�yX�t�z�+��>�D�N�:a<�]ג\���m���U��\�ȑv7á&��DGH��h��Ֆ����p|��Oʢ������n;3�P��\�;��2���}���6:ְF*��TճQ'R�Ǘ�T�̉F�ɘ�zPYߠq�b��`s6������Fи�����/|�A�Z��U>�s�\���ż��������)@���8v�r]���'��7�r�SWh��L����G�#�'a҇
QE�P*�wı�D;()KB�{f�S��¢�^��L�?Z+q�X�X���c�<����>���͋��7_w��_��V�^i54Vr*u�ow�g����~���y���˦)�@?�e��{������b��ɢ��p�ʅ!��S��#���ظ��x�����v�?|�P~��2Q���?�8͙�e�LچG��g����M��K��ƍW��;<�R��U��̳OM�8	:l��z�>�5���w*�_�4k��K읿�v��l�T�a}G{o�J�d�Lڵ���CL[�i�������y\ D� �4
�cҵQ �"I����w���hf����<9筷�;u�ی��H���;`8���q`�[�Ɩ/���|�����7��K^k��y]�	�Xiˊ�bnЖѬ���7�D�G;&��_ו������	�����?����^����-�ͺ����l��:d��r\�[
�h�0��A(.c�x@|�3���'����J
��p��1�x������c	��@���IL�
�M���� ?�O�u�[V��T3���<q�>���5sI%�Z��nW��F/�ݺuvͳ��|�l���dl%��C�8ξ��x~���?��I����eng��f�XC�x�T@ɲc~8�d�ŋ8M{��I{��'m�L��ǜV�g۬X�x�E�����l��%�\����V�Xa�Q�X���i�={�xhh�����dO|��׿��v�O]���~;u�=�k�ϟ�S'�˲�H�ldp���Z笥����c�S�cO��dN���N1�_~4�OZ���:�)�3���#g-�L[&�a==��U��86��&������ݏ-�Ϙ@��1�R��B�㌖̢��������LlEca��b9��7{��; �X�YE-���͋�G��x�?�2�gh�>�`��gº����7���;o������ODٽ�i�7k�����)18�y^����ONe'#9�6 �� �!G�
����B�`)�
�F� ��/��K��M��ۮ�-�iX�D+G�ի7ؚ��Xjxm�l6�a�����yFm���(l�&Nw��F�}"m��G졇�^����J@맪't��uyn�
�U�kTG��w�����J�UR�V-��[�a6^(��c�v����7���$��_��_��u�Ȣf�'.�v�����/6��O|���=�������&����Ä��}���|�b�U��o��/m붫lt����?�ٰ,5AJ劝<~ʆF+6p�lo��o�9@�Z99O�c�������R�?��Y�<f�d�Μ9b�=k��l��Y��?mc�����������㣈*7���`��%rg��s P6'��E3f�J�D��QCu�K��ht<�?�g���#��2��ٖ�[=�h�O�s��#��ޫp�2��١c�����J�'|O��BOhМ�c�	*JH�� @IF���}�"@H�C  ����]@(@��	T��8��|��O*Y��������K�Imݚ�m���,���*�`=_B8�;:]��5�8|Q* ��z�(��o}���X;U�|G()��k��<��J���=k�ʈ5�e�;�g��H,sK2�fǏ��b�aǎ�[��N۾�j��=��<H�G��d�ό�[���������J��{����ۿ�V�n�j�?�h�]���"���b1r �r����<6`��,;|d�6l��)Z%� ڀI��Y3�ACCӜULG��^�÷2^���\�a=={���V#q(�m��� �i�B�2�>�l��e�F�9��h�܌;>8ru�b���,B�(@���d�Q=�lp�)�+ |��;��/��"��=�:B�G����@�a]P3�?4�# �5Ƚ h-B1�.��8�cD9�
e��\�*�rh�q�����p�N���`9p}�'h�XXD�`A�(�(i��fM��B����i��E�D����\�m�Ԯ޵���%��m�u�Zd�_q�Y��J���HeL��'�X�Fl|�>���@1����o���Zd��Ԕ"� _!����c8~h�����l�ڥN=��+ǭ���}
�Z���=쾉ѱ��Z�����wXG�l;yj��z��S��[v�ghx�C�4Қ�+�W?�^/��ݳ���7��y�c�{�4N(5M�mhpغ�{�����c[�&�I�X���h�T=#��DLl68q�ԅ<�ٜ���p���IT=sq�8lgN���[+�[ �筯�k�����sV_ �_�3o��4'8{���Q�)�q%�B�=�*����P. ��������誉
�g� ��C�q�j�ε8O�;�& .JJ�E�9�/�%�&��r�u��T�kI �x�St���C�����uT��5۸����|3��KY�e\�#
�$,a�PO�8��������_*[.�r�/��յҮܴ�2�v��	�C@5��8~|rQ����sv�0A�1��94|�֔2���r�X "ð��������|�6o�`����w����b���B�n�=w�2��v��/7�S�|�
��7R����۩��x����u�݃�C�>��=�6�j����T�f���}��u����^�����6>Vp��d�l���9r�R�Y����bӎ	�gS�� W����H�4�8�S�Ntc�l�yq����D�j'���=�X�FB���Ȓ = ���z���J���X�("�y15-�8z��[�x�d2���_߻�4Τ�,��TV�����k�������Щ�s���y�����M��Rք�		��1���ֈ�wx|�<�YϦ���u�q�[���Tb�����*߅��`_�g:���/Xow�����l��Wx��<�u������k�o���h�r۵�Z��Ky�Wwx{;Ԇ�������D� ������U�ư�H�D��̄�B��88�}��_�(�9sf��C�}L�wTm߾nK����Q+V������jG�#�K�qԺ����En���}�|bhh�7��=&���������w��_����~�N8}�J�b�O��P,ّ��66^���5��ҫܳ���I6�q��MQl/�+���(,���*��'~�^�h��>���O=lgΞ�������:M�H[6�n}GO۷�����,��l���d�ǛX\<�o3� (�T���&i��p	����څ]\"A�^��N�y�ֵqB�-v�K�I�&���h�uX��.V�tr��}	E�85F�v���,l���8��^=ח�YA�r��zg:p��y���m�%�b���'�k���C͈���ވ���uA���n	+Z�Z�(�T��͌U�)�5�~��W[��o�6+�	���x\����#�4�^4���}L�oYc8�J×D>�|'�D�#�����)����b��-����?y̪��[��2/�O&�e�N���K���?d��s���1�����+�_�p��fjI����gQΞ�i�|��l��%�ޖ���_�+�Z�6�_L?�;��Œ�����Ƭ�t����w�㌍I�6&E����LD �S�� ���jT�W+��h�,sm�<qB�9`'Ou��\)xUO�Rx/��}z�>i��,7:�f�r��?tBJR���M���P|����Pb!�zC�V@h;��&�^Cm\�ǉ+�Ix~��f�s��4��u�P#��s����9�/IJ���P�,�����	�PP��-�f�L�j(�4�\;l��K��b��Y�{����3~��8�{����|.e�zɮ�b��ܹ�s`���wȵ�{M���k	[�z�U=�&�}/��I|��>g��/����;��N{�k~ƅyDt1O�����N��O��r�>��}�ha��S	;5pʊ�1�1� �z����q������7~�k](}��G=˻T�|�/��$���w����Ї'���j%�F�[n�����6V�F�h���sV��G!X4s��e��6tn�N��5Kvٛ�����<B�T��E ȓ~Ы�
�:�Y({���I$B�	gQ���*�P��>Lzil�Ν;c�:����Y:8�̒�W��И������k����k�y�8�E�}BS?����� �ٔ5GY��k~*�����E�7�����e�:�����t�/KA>	���-�
QNa$����)ԶC�Z,�@W���JX{du�,�4���JP7[*/U�!�/��kVZ�&�?��7��O9�R�9]Y�;���uG�xT�����Ȗ�x�t�KĹ�X |::���@�D��������O��!��R����������ر�����;2|�
�v�d���7Jʹ��:�y�IK����s{�E�?�V[�d������w����po�
b�^�ɝ�n�����M	���Ă^�|���]�b�ͷbaԆG��#�|����D#2)�eʽ���c��̳k����L2�rl Ջ�!�VzQ�S<p�lZ8B��r�h���6�&����5��g��=K'1�Փ��|QS�0�k��B�H�Y�v�z3��	���"!.�� ���7���4�f�#&ː��<iѡ�>ḇ�G ;-���}�Ly����.��9�C/C�<�eB���Ofq�<�q�Ӹ���BJ(����T�<%��f�n�g�Q�����-�({�Wi|��u5�Q�e"��b�b�sl��^�'s���p$����V-����)��p�b1�Z���C6:%�(#��(!�����[�*6p��>t�N�������6K4�^_��Jf슍[l��U^���@�,�p�M6v�Fc��h�x��TEB\�u�ַ���Fm��.;sf���N�BR�}�Nۺ}�D��K�B���u�?� p|�m���P/��<0�	�ęL($Rǽ�b*��'�}�8���Þ^�j�ly��b��6^�������M ��������{��Es�����oH?4[�=�/� i�D�6-�?3QP:Oc��!@���|�eYH��y�V��]�#��� Y�u��K��*,�&�3�4����v+������m����L����E�H@�X����,YBmh��F��XH�@�.��a����z�T��W�	��I�ܰ�J��[�yKPJ�����w�    IDATa�1�>0p�>��>g�Ҹ+R�Qf�*�K�w%��P���	�ݳ�+�
֖�X__�=���=4���âF�+V���o���̙��B�9��E9tz��gF��n������_�J�WU�Z��Y,�{ӊ��Fn���I;E�0o�Y���p����=���Q�(&���:���P%,TZ�7����T��@�ؖ���5m6ɲ 8@ǿ�~�N��X��=q{:�p���{���=f�c��f�^%��[�bu$$�+�x�>���GH��+c�����;�R���m�N%<D{|��K���t/Γ�PXg���<��s��9�<r�N��J
�yo�y�B���C��g���ZD )�?�~B�*O�
?�'�����][�P��7P��J�D��U��j�T#�?����Ջ�}�e��͖�G�I���w(������1��"�oo���>h�����y�����w� ����16�C�w�hb?��
7V�U��`���J�IgG�G���%'%0%�����xN�9h�o~���v,��%�Qѹ�>3�o�s���{%�D����.�ȭ[7{���~����{z�%HĿ>���.��nB�S-5�&,�E� `A�!J�Ϳ{��y�E�ڏ��T~tޟ�rq@�U���,۾��@�/�z�liZ?&���s��i���R�膜7���K�)�-.nIg9 
9cƀM�u���D?1��Y�*Q�xJ �2��/ R�fb��p"��P�G`c�q<�AT�^c����9��p׆� #ƞg&v���]�~d��X(�D�l5�x�,lz	M6� �g�W�%����[��{�X��D�����pMţ��Y��	���?W���M%
��g,�G�J��%ͼqnX�q$�AIz/]������	O�"ڇz��,А�y^}�&+Ǽ��$v5��'i�5{�]�e�G Q�n^hހ?-�3������w���ٟ?��M���\@��G���}����Ԍ��E����[}	%oԫ�k˻J��7�I%��D}��oG�qw�tTl���,����i��1������+lێ�v�����Ʉ�g�r`ч�t���A�%ٚ$uQ3���L���OD��6��#����[5s����#�m�T��k%��F-���B Q���}}�v���c�굤�]�>���{�.�CI[�j1�� �f �qz!`�v�V$)������a���G13	U�Yuo(�FF%�qŜ�: !ay��l<
�~+͘��l	��������͍�M���4�H ��zTڤ\��}�A�l\(��F.�$�OB��|��'�G�Y�Ō�Z6�.܃�PuX�EX�=nٲş�h
"@�*V$�+�'������Qh��'�źe�B?��Bk�8� Y`<Ϗ��5�j��U�P�0�{'�����&�.��	���Q=���m��N����^�皫7��)ژNd�TnX�m���3w�OC��:��6��j�Q����g����w�����n��V��#ܓcM�?B����߉R�>q�w���Q�Q@j'��")���ɧ��y@�Jd��]��'��L�󟺼CӨi@e�+CVC�c1���dܵxMJ=������I�' P��?�A��{|)S� �0Z�����j���9}�z?g�҈�57sm]v��xTۇ�΀������3/ry�K���j	���Q@���#��	�c��ËEŘQs���%@�	� 4(�����E�y��G�MŘ�`G���G  Ҙ�gxX
�Q����� U�m�|��ا?�ihr4e">���fF � P9���F+$������^]��C  Y�J�`� ̈�WD�.��@E��]��A�I,�Y#�1`iV����r8l��y#f��C�I�����Ġ&e#�;�G�ERm���<�04ɅX-���� ��$�"��*��9����g��zz[6ٰjm̶m��v��̊��FK-a�L���Zn�6l��IZ��Jw�jO�?<;�V�
��}�3 P1o{���C�kpg<QX(�G�&(�ЂcND)�*7�NtR@O�'�1�¨�h��o�u�g���?�#Gd���Z��u՛9_E�4K_-��-@`�g�e��� h��[����W�j�d]�.��������iTk^ҹ��ɉ�nQ3�FT������.3� '�ECcs��Y��� �G?�Q{�k^��-��L�� F�B[D@0/l@�z��Z�	Z�� 	@��Jm ��4rd����c4��kM�b�U���<� �l� �(�v-.B:g>@(����;k�͏@C�N�0@���Z@�G���'
�!T~4��ތ-��&H��d]!����ð`X�|�*���I_c��cҌ	sûBePH��5<7�KDy��"4��v�!�0@h�>܏�X�|Tj�#'���J:������@TϿ��r)�re�vn�ܶo��C����<.���XǬ�6>^�j\ٓ`	�ѕ�j9�ԫ^6����
���}�{<��g�b	a��֩�
�KM	X�5s�5��q�~���w�5�x�}Z,�j���XͿeU�x�B���P (��9�Z1�!'�̿q�����j���aΫQ�%�ܻ�����e��O����Nؓ������rVk�����#66vk��bY�����{�}������VҏLd�l��y�&
�r���D��� � ���1��$�Q�8x�cs"\��;�U?y>,1�h�9�ȓ���Ei�*;V����$n\��h� *-3P�� k �x���������]w�����@�g=�BQ	"@��L�6M�i����]ԑ�5� f���tPj\���E�	���L l�������a�b��bC��@�1N���xƇ���ȉ�����'̎n�W�6О]�$�����L\�?�ߊ����k��+��}�Wk�^j+�\i�:%*���4�N����LD�`&�t�A<V(x�^��GuPذ:��+S�RZ{�#��X(B4��/֏�����G2�5�[v�~Q�\����hIi�k���P�H�7��\
�G��;�1�, ���%��l��ג�M�^AC�ٹ���'�F�>�ԸOؑ�1��MN3��zRҙ���3�p����d��w��0XGP2l*U�d�Uvm ��PѪ��DB�;>|  ;�8�0�k3)���C@��riV�g��M-M�gCp��w�s�� �?��s"��]3��n���~Ο��������D���Y�\��P\��<��E�@��z��"� ��yg���̀���JQG_,,31��5�c�b�7��1�Z���`e�<ļ3�h�X#<��1Y9��J�\ɩ�B���������|�T;�k�F۾�rK����9��z�[��*�6�V�'�A��Z�����#~�<�b���r�|�9ғ���wG�S_|ƞ�fܨ.���|�~��0�K�-�I��!� ��hi����o1N����wF�����#��T!�#�r���Q6���ߘI�\hQ*��h��X
��h���k��7,�6;kǎ����yR�s����3�?�����������F� � ��)9 d��!�D�������C�x @�#xo��c��E�b̠'�ș b +� ;ԉ����� XC�\_�	�q�H�h68���������@��9~�"���t܃ka)��o�[����g�Fk�Fh��:2�� �j��
Nj��x���NW�AG��}�N�O�ϸpm			F���X.�(��@���c2�|x&(N,+Q��������&�d*Z�����q��1���*�^<����F�*6�R[�f�͞���;$29KT�zD�e,��ɦ]������>_�zT���c��T�9U�g�{	נhq�a��K�F0�\Kʢ"�Z�����n���}n�whh�=Sq�tih��Zf��t�Ĥ9M5��|Y ���hB�)'����A��7��ꓨZ�6j��!;s昝8�cV�!�_	�Kz��Ѩ���>4��G������@�KfY; �$�V\04`�JX�M7��9�GÇfPC�8�~E��^6��0�8�c�9�s�����8D���<#߳�)ԇ6�?�v��X�Zͩ�	x�ݰj��p�h�8����K�X��@ A�`=�}�4d=���7�e�@s�R �yg�1��yXT�3�$~���&4 ŸBc��2�9��	�*����!|��4R�C� �emx�z��~48q����2�p✃pVn��k̉O�S���9��Ba7���{���Q+�V����d�ƸY��c�,a��$;q��<���ͷy�;��h�T����;�z�h���P*<4�ֻ��Q�G�:o�@	;�£C�AX���J9l43W�e����{*�,���w�Tܿ��Pp��C�˹����5YD���s4$L~�^���0KT���G�T�eSu��j�&���NB=�����oT�?k��<� ������4PQ5
d18E����� Z'�1c�E�3�aB�) 8R����	x"Դ]4���
d���V���������w<�V�/4�k��b�p=��`m�vۻ��?BI B�{Q����Hy�6c�?�*�8[�l�J��G0����;����F���?A�T���gM3X<�/��cqM���r,ϧh"�Hh�r�ù�0h$�3��
���'��O3��[OOTҹn�y�Z����I��`Z&=�GJ6g�����a)��I���l��g\	#��λ��9ͷS!7:��yY�
"�~������؇�������l���-Xxیl�8�K�ntw�0�q�prB�j�2Y^2��[��8�l<b���h�o�bO?y�x�?qι4�a�nƶ��0���o����ڻl�P����g)�����S	.Z�DHP�Q22��R�o���3����^�"���dI�����cj-M��C�h��+sqmy9�B�D@������~���uq�P*PC�,��D!�y��XD� ����=Ѥ�%ᫌ�Ve�� �;��b�f�xVU��$r=��wFH��ܛkb0g֢��/���a�w#��5˹ⶹ&τ��傠��X��"��S!C���/њ��D�Oe��/Xo�a��?:v֮�z���S�l�0�;�L֪��n�:V�,���WY*M[Ժ��qͭ{�{��G�c��Oi��eh���B!�5�R�C�����R_g�
��֘07��ߕ��
[�y+����U`�s��ܥ}6[�'��,*�k��Z��1���N����A� �w����W-Q/��fuം�,�b%K1��ځ���Ǟ����'}���r����b5s�F�C�$�Yc	8C�����@���Q�ތ!�E�	�7��ax�"M�0И���$ņ|� ж�x�T�.�A̛�6�^f;@Z#<a|j̃���%�Z� �ϵe١y�
�û���������]є��.PK\ޝwCx�[ ��&?m+�֋�5�D�qo�K�1�r@h��:NYuSh��W�.�$j�ga�3P]�{��	�����Ԯ����=�MĚ�y�5� Z�w�*��^�vݼ�&8��+⪞�"9|)��qGj���M�m��+,��z�o�ޒtK���Za�dU/�\�|[�;~=�2���pl�+|��&ٓ<���\�Q�F�	�sQcr��]�5\g���p�$E�_�F�Z���,\����җ��������i��3�,X����Z�)TO&1�b�i*�xX��X��o�y�%幷��l��Bi6�j���h��IFo٪%
WQ�6�`_�elp�`�D�ʕ�,q�˗-�����0�a.tލ�6?!��s -�b��@	`@q��Frt�'����� T�7 e�����+�G<`�#�EH	\4�2�����hL9^��O���1�z�C[���%�U���yމw D�l~�#�����>Pp�D��`�6M�)`������P.��揟 ��Z�̬]�%|%aƅq@�p<�
M�{a����0��<B�s�P�^�R���A�u�_~Q'-@��\<�g�
/�|��D��Mٓ��kE��H��Ymf����)����@�'V�&��HY���\�͊�(@�8>�}F%�P�%ӕ����(2֒
���Pȅ�(�kM��0��f�*��Y����o��o�����ӄzJ"��*�]��f`s�  �]Z�jvȡ�w �4���S�!�P�tp�:F�)a�`���CV),�m�yu�(EͿTI�h�j����3:-_F���.nw9
%д	xW���`C! T�5 ��ln~'�@�)��#��i�r�|4t�08�*<6�~� x.�A~��&����>D�i��W+B-\�7�E�p}�(izh��MJ�뉱A;�U�F�O<�:�j�+34
�B!��/��%�9Z������� 0��DQpO��\0'�cM2����X�#Qb��S~"�p8�ySY
���r�<>#�V Z��h.�d� �~X4��XOO�u�wX�4b�d��U�4<J[��h���g�Ξ��6n�f	�zE���1��eU/��"n�駟}��|ܰڇg�0�����1d����h3�Z�̍���a����1dO�\�l�߳珇�o���+�����ĝ�Q�d^n�^���t%"�́F��l��
ȧ�Ρ���-\2��*ɋ�'��������Z��Z�D լAU�l����g��R#�n�/Yk+�/���HR��q�Ffч�Ei��5#�_��4om
EN��F����Fi�:�ߡ(�#E\pOi[�V�����

-/��d��y|�dѦ���ϵ���s�4QMat����QD��$�Bk��d���T�A��,S���hL�!ϫ,w���3+��Q��9��q_�%��k��Ƶ5��;O�o.�����cL�8�S���s˹�(چu���K�X�:�e��(y��i��;��x�n�V�}��N_�"h�h|3n�}�'#|h4\@Wc+k�C��;�
�C9\�1W=)�%�f�0D`C���A("4�(7~�20�OD{
���Ok���f0����%����:�� *�y4=8LņK L�
56�xa��{�c!���I&jv��S6����esIKԫ��ʣ-:���}灇md���x������5��bT�x்.��ؠŰ��=���yKi�l,�IZNH�79w%�Gi�y���X���ϩ�' �Uǵ��#%ABBڜ�Eq�l��tM"kI� DJ�~���7O���Z���9�g���y<oi��IWֹ�+t�A�r@r��Y'��X1ךC�'Q������ʟZ�Mt��:]�l&a�ڸ��v��tnT"���m�7��-�=�����:w�9��Yq�lt�i�Ko��;~�-���7�4AI���� 1���"k�c�
&V"V��=QG�&(�'(B�>�Kx%`*v�e�o��3	�+76��8��Xf��&4�"M�c�˄�z��8��H��{Q"'ؼd�NI�$��w�#6<|��U4\VQ�p����a����~�
cKg��J8��{��b���N�"�i�r�3C8��j৸T��j�(|�kl�fB�I�� �����p=6����k���mq���G�&��E �@��8_Z��$��>�X��:N�������B@E��}��r_{�IK0!Ƞĸ�4x����(���}=C(�$����$���CKq* �{Pҹ^����aˤ���!�r�z۹�*K6"��)�\�P��l��e�e�.+V�6,��{�&���F�-�?���>h���֬��N�=e������C �J�#c�>Ƿ���^�Z��QLQ4�����/�����>��>�B�>7���v㍯�&<I)�aw>���޼����_h[�l��wy��5�IDy`�� e*����A��c( �*ԓ�t�3v��a;}����/    IDATU�c���(���\~����?e�Σ�Б)�&��K�{}.V��(i���%8F��%zi�i��t!�0�3��K�4���e���I[�!(�u�*�%���s�kB�c�f,����OBCt����9*�gܸ�'�{*��"ǤK��K )�M�U�c��)�� ��Ѹs=	EJ5BY`�B~ 	E�I��&�?/ ������D�oV�M�а7Z&E�fT\.��]�,�d�lպKl���f��&b��'
�������OM�d(�K��d,�ې�Cd��Y��ɾｷ[[[��mY/�|��q{�{߷����o`Ū��;���a�t���Pw�����o�/h�/�����S��K�w���p�l�D�������Ν0h��� �U��⥫�k^i��Q�)�q�L��~E���ӂ���Q{<9�ظ�>��V��&�����f�L�Ϟ�Ç��b��k�C�g+9v���S���;ԓI^5����o^��¢;H��Zn��n|��@Z&?�'p�w�G�d�:�j����- ����F`���l��d�9N���Ӑ��=��7�D\O�o��hQ$�^xvmx	{i�>F��k~�ֈ�AE�	h$T[�~j���� ��.�z&���%�{zڧT�m[/��;6y���r�b�d�.{�.�5w�e3m��ztl�#���z�j5��l�C���Oz�s�LFY�a���5�ߎ+B]�Xw�2BUٕ+�Y�R�Ju�~���l���V��-�H�u��>�.�|�m�~��)A�L�����O#k�g �V��=����F�x	�¼��֭o��
�C66|�N���޽6Vt�ϻ��='�v����+I�;o����q��r�<�f$�[���Ą��O#
ca�
 Ĉ��*�� �Q:e����ؑ笧�+���\&c�|�uw������6�sA& ��F�L�A�����H��}fuF��DE���V�(c#�(cE�	ILQ��W�6E8'@U�i��[�7	ݛ���*��n���s ��Һe��9
r�[�{Y���k&�ώӏ1����y�$넱iV�uC��z���Um�����q�'r���m���M��b�F�/]mk.�ʒ�v+V�^�'�J{/���X�)K�纎2��Iu|�Ɍ;g�KE��z�����{���g���;�����ș�G��{�<�φG�hR��
R���F+���]��M��	+���hѾ�կ{QH��~�VY�/gny��J:k�9O�_�h���i��?��-Y:���<u��e4����ㅪ=�o��������.�p���夝J��-��c��6�8T�>$<v-7w#m�T�����Hة�����,����$g�ݪ��&x~a7�FKs�����'~��S*VX��ЎD��8�\T�����U�� watl������Bg��q�lB2Y	uĤ�C$���$�!JK�ҶC��{`��k���;D�8%�qo���x��Y�8p��O�h�ٯL�� �N�	��O���d.�?Ɓ�2j"ϼ�S�p�a��/O�U�|�R�Nh�����?��zy��;7Z>mV$,�Ҷ᲍�pɥ��tZ�R��D�9���9���s�t2�@Nm'������=���y�X(z	�H��LrY���?�����z�F�O��O���Ҹ;���Kh����6pf�j������b��^����}��H�iB�_�I�t�\�of�aK/�z%��R���'v�+��$M�{�[�i����cG��V����C�e�.O>Bsd�PGF&�f�_��8[4?�<�Wm�B��>��U+	�fR�˖���C���I�T�L۱���f./,��O���0�����O ��fc�H�v-���������C����p�#:I �Xq��0����>e�)����x^�&d]s�� �ʼV�l�"2b���z>6*N8������%�9aA"�W6̝�"	LDl��u��I��Z��#��x���A[�j�+!X'T�Ĺ��#������Ci�G4�L�LK����C3�-�.�]�l�|�zѬZ��K����vX:�?8��Rz��>$|�͒Q ��4��mDh�];=�\�H�#Ɏ5E2�Ah������.��w����_�����C����s>�POc����{�::�ّ��v�ƭ�����^��pw����:u©ח5�Iv�-{��l�X�W<Bf�ʕ�[��[�j��ࡽ��w��j�g�8��&�D=i�#E;q���>=G���;<}���Ԣ�
�(��d����pO��� A{�yal-�z��&��l�'{��@��=s܋Y	Eu�W�OU����1���S�S��r˥���Xp���h9�È�j6象<���pp��.�(�' ��LZ���'��0��"��|
��tE�.��JHK�秢v�`��D5���`�����/x6�9��<6w��-A��P�L��\_���A����~e"�MO$��:�*�#~r�>ƃ���ь�������j�yrc\Փ6�1��s	��kǕv�5��j��UzZ����m��E���T�?�ō[-f#'>%! tJ�D4e5Ŝ��F�&un#󙪬R�Kb�c��.�?5��Wl��ˬ���{�.���3Y2���S,�j��g�-����;u��M�pj���!�
�̥}��d�F�%[�z�}���3�(��O����W_����w�5��d"c�C;v�U*i�>�?Z��o��J��|���J3FC����/�뿣ɲ��rQw��k�^.���3���g���&�!��N�[w�@Tҹ���Z�Z�}�����Lg"39t���+����dI�h�	GlowNt��elr�)�S� L�LS�js��M��B�@��	L������|<;N;@\8s��]Ř�;����u�������Z|8��9�g���|hͷB?�t��Vu=5�x'��8`��6

�$�D� "N���-���pή��*۱s���-���IZ��0Kϲ��V���Kl����9&��F"�0S	s�k4�.ؙk����	س~Y��]��Z�R@�,��s���y���X.��cǎ����HФ�ܡ�G����ђ}��`���V��Mh���
��8c�8NG��,��d�:�������u��/~���~��2;ܽ��Q�=��C�#v��	�V3�w|Զn��5 �^�E#'��@���h������{7'�ςB�g���� ��M�$��lh�%%�g^��z$��������X�Ƒ�nk��ˋ����
� J}�G�$�86�\��X8/��:G�XDu�0�Rܚ���<�� :�%���c<�7?
J�P��&��͇&L������A�����q��=T���/D8V��!U'+�9���ޔ��܇�D$�p9�~Rl�|#����(�-�$�Ph���z��Λ�q�;
��}�9��7�у��
�]�H��
��$jhZڇ�==n��#v��+lێ+�Ny�l5/�l�U�d���]`۶�Z�J�9�T�lg�J���|��]wOXz�e�4��p��)�֨ΊR��l�)|Sp�(}}{��o�/��ʵ.zz��Z�!�����Xɞ}%`����Y���5��5�N��v������T�`����f.�3|�!��-g����ys�X�������֯_i�cC6<�OF�����;f����l�n~ÿuPB�S
�pO@�C��P,V��͌_Gi�L.jD.���E��M�qPKT���'�H�~k�S�d�3}]�E�I�[O7���9�����Y��<_��W-�kw�zʣi�_�-Y��n�G&Q|7��MC���p���h'~2n}��@��]�M!�F�6 ,�	�Bgr�+�J4WsC.�6s#*Fs�d(9�$�(d��z:j���J��C�b�K����8yk���߻��.�8ʹ�����.�}>@��%��`�'�7�}��1��_�mۖKm�+<�'A�;B=3yk��l�P�9�ث^�+)~����~b�� ��wMT��C2( ��)�>�$��K��`�}�"a�(
��=��7��3ms�̲��38m��y���#�ldt��O���ڛ�g^{�7�yv�>/��E,+�e�o�
�U�L��J���M7��n���f��k�#�$h�,K�?[�9WΟ�S�m���������S>�Z`�q�UE8A�
y9���'��aѱ8�j[��U+E�7��P�8bV/Fez)��ى���s�mx��>�锭\�ܖ-_9�����_�� ��r�~�~�ߏŷ|�R���W��Lԯ��"�І� �z~�w~�#��}����&���f�`m�	�6�h� +?Q>h�,|��\���&��1/8e��XlR����1�jnx6Υ.��k hb|$4$,ࢱ��D��I��d��q�a����PH�Ї�}�O�����w�r5xq+%Vx?�k��1�k�߈�Q<7�w�>����V�h�t�๰4�o���PP�;���M�>�a�C�#Ը?����Z
��x�� ʵ'�L�v���lTҙz�����_��.�b�7=�륚�sY+��R���ZmX�FV��Q �RX8��t
�>N�5���N�@7���ظ+����cL3醝���s'm��Y�JH������1��=f#�{ǯ���`����}��}Oa�Lc�-X��/���|�L��9u'�F�J�Zd��Kv���/���6����s��SO��J�FTK"E�� �,�]���;V�dTT���Z�1�p���lf���" �=�7��b8�y�RqI�L1���U\@5j�*{�?B�\%3��,w����96^"d�b��|��X��
�޴���}b�R�ģ~�	���t�Zf��t����h��i�X�� �u����ȣ�� (m@J��!c��� 8����В�3�X���&��y�&>;Pо8_t�TH�iL��9<#�}�K_�,����0f�a9`��� �`��B@vZ.�l��=�Ԧ�	�L	`ʈ`Ma8��J�v��: J�φ�2�D�!�yg������.X���˚�3�Y�Șk��z�|x�3���5��FR��Nh#��yg�@�E��q
�yE��T�a�^��d����d�$�����V�|J2ac�g-�M[��4��z"��(K��-�J�*�/{�$<q��dv��T����xG�Sy:�8S�R�(41�˹0d�iPT��[W{�|�z���(�uKeӖMe�\%���i۸y��[{�c4�_�K�7���Tz��;s�����}ph�]2��xs��HZ%n�<>:�����z{���R������������������a�V��׾�&K��zł����U'���bƹ�4���'N�t�s�� :6��<�q�8M��mu�?q܎�v�?�%��:��L��600l�t���B�
��X��J��:c+�'��;�t$!pQ�����fuL4� \٬$_1ԭ��"d�D��%2�1@�ط�9S(>*��;0�h4"���k<_���ƕ1Ҹ�a��3��x�d��0[��b�)�E�C��*j&`I�c�I`�d/4Hx`@��[h�p�1T�7���������h��8����XB����.�hu�s�?����ܯ",5y8�G��p-|Mh�{� `�����u m�lƁ�&8l� jd4Z�\�5�����>��D�0F��%P憹b-  ����IP������V}��k�9s;�R������V'E��t�=�6o�f�k�v�Xs)��	�60?�G>�)�(�x�b����%HY袁yO�x�޵Ò����{�g�'�ǎۙsg<�c��Ev٥���l��n��Dʾ�������}��E=^�IF`:����|AΛ=+���|s]w�5�������>�4�����uk-QoX�3~�644�?4�o��f��h�y�r�ı���h"^����ب��	��ھ瞴3T�L�,��Y�R�Q���t��C'�������^��s�-[���5#��Bm������,b�n"�`D''�l��e3�b����Ip��Izcs#h ����3O=�&36r��9��	P#�µxv	�x������2��46-V
�E�/Z4��D�V�GQ�G�]�[�/�����y��Ra�� �x���&ƀ����# T�z�k@��X^��>�4��LX_<'�������1h����'?� @#��C�@� �8�Ʉv��������Zg�c�Ag�8?� gm�[�_��`�P��(@�o|��'�SZE�fj����P��>�4���2|�N�@��֟���x��/Xb7��j#i��:���eg|[<t&���½h�B�19�qd3��#ㄦ��\'�(w�wݾu��!��(<pp�����  W�Zg�]�622f�]�큇h��W~�H�L�3��۪�{�0�h"Ж	�$������WU�^6��ѱ1���v���kAl��,Jܒ��F�q|��؀���������`)@�xDJKͿb��>j���d��5~*�B��l��=���=aC�t����YV����ޭ48����Dҙ��>���'lvx�
`ġ���O�k_�:s���׿�5��W^���F������.n���ccqc(�l,
�b�� ���>�FT�]���VZ/�B�)�/�e�h]���Q��SҘ�8t?~z</c�,nE��,<?�����C <�ll| Dƒ{2�h��?����k ё�aJ��̀P�3�!<?���&c�u��6�;� J����F9��`y�����8Xdj􂠅��:P�Xm����{� ?]�L������"�Zh���t_j_U��^����Y&I^J�Ն%3Y�d�FƊ6{�|���<0�.x(:XfШ�?�K��p_�v�ڭ�[@�yG��S�>���������׽��8j���A��j7�(a�"s�\�H��������w��Q$*�MHw�O��(�\🦍#`Ƅ���h���h�L�Wl�-���Ƥ�_D�@E� �*�M���j`�"�p�hЄ=)a���Xm~�v��ΗҎqJڧbGz���'���4�Q�!w�&��p�){��O��%�;�Z��V�p�GV�T�?�@ |�cI{g��n�J���=������G�,Z;|�-������Zԓ�?1�)��q��c P�u@T%m�t�����"���wm8�ņ��A�0�r��@��.aYO�<��q�D�@�BQ>ʁ�'�O�K�s \z�AK���|���s�m���#��oG��G�=���Z�ǃ����f�l�a��5�X�PwX�� �h���g�0( �\���u�څ�йV�� �=��P�Ϛ�jb,v��I�'��xX>Z��͍����f��;��{�r٤U��z�z۱k�%�eW�Ru =m�ɜG�\�y�ժIKeڼZ�C����G���}��_�E��G>2��b|�g,w���*ժ��,T栽c�]q�+�b^�v��x��G�`V�Ç{���r
S��N�
��gl��t�>��,2@�	Ne��F�*e�1Z8v���j�}#��бǩK��Y���9j "�z�$XR��?Q�BB%�[q����lxp�FGO���i�}(E��s�Ġ}�[߷ᡒ�ۢ"j ��UK]�F�i��cݐ�Ef#-���/~8e�Xo_�or4B4M VM�т�� 6���骫� �	�-	m<�m��;(��h�|�8��8��^e���f���]������N�7�6�W%P��`g�a�+GA�E�T\�(#9|�;�׀��g�~�%�)*��b�������}��|:
c	��Ppli<*�O
��u�������r����sq_���ZQ�@�J���zrT+(��eMqM��g�r��8^TG���O��Zͽ~j>� ��)3|[��v�����
۱sS��e\#�?a]]�mΜ%��5�/Yn�z����?�L�ӗ+��>�G���E@~�w����)J C�bY����)6R��1    IDAT�gfnU�;��f�%B�#b�����K/qg��X��A7��SKD��{ǭWy&/:���?s���;��/Ȓ����'���ظ�e�У�^�s/��p
K)Ւ4���b6�������ܤ~�m��T��tf!Q�`J�oDF_[&�)�=m�O1_'���#>n?�d��H[�T�K.Ygk�E叧4�X�{ m���F�n�3.�0��~�X�[Ex�A�Y�߷ϳzh9,l�� F@���G����E�1D}��|������A�I!P,a�Q	�ph> j�N,5Ȁ�����>����.�ڝ|xfq���tM����a�����W�ʩ-��+?s� exVh�2��zr����"����uO�����&|P�z��»�""�k=N����h}��� <�ƃ}��%�����; ��<�s4��/^Ѥ���h���)+m˖vݵ���;!��x�ƆKw��+�^��;��A���{�tųR܍����r�{��`3� (���r�χ��KOF9@h��e�q~'�8B���3I�����"��C��7�֚d�f.��t�Ʋ4�x�ġ�?��g�b�4C���D9hCiSPd�@5@6/+��s�펅%z�Ο�:U��H#JZ:��.^�D���{��g��+Ke�Xo�I{��ld���Od@�l�b��}����X;:�"!��c����B��[�0�<!nJ�
5}Ox�{Ȇ�����������T�V�-����t�{7PÇ�P����59_�V������\�MO�)`h*��s��
 6�j&XQE����_�U6�m��6��::8Xq,����/��}�����d��<q�>��(×���d�9j�� )�IYq�d�/��V��l�R�uJ_e����q�6I�����]�=Y3�j$0���Q9q4�tsnTc���3��?O��1g�k�{p��-{n�����`���y�����y�'6������U(  ������
����� ��V��  	N��h��4�G�U[.e4j:v�:�Uk�3���}���>j#cD-D%�q��\N8be��Sq����.���=����*m�����݉R�g����N��V�2^i���xL N�WtL�M�gCX�D_ hy �)�ĵp�J���j� /Z8<59��f���¢t\_�S?��'���%�-����Z 2
��jG7�waX_3�s���]iU
�ў1�
��ϛ����q�Į�f�%K%jV+���ˮ���7Z�Ay��[���(�V�|�#8{�O�O�uwT�5��=���DAE&)���Y?-�gk#0�YPJG���r|�N���Kj���{�ǳ��<ON硝�x ��O@��������ln�"�Z/덨�U˦y��uz�z�z/�l�͝�ǎ���<�Hk��zfŲ�����2�3n�ieq�}�t ��C/8��Ǌ��Xw�j���CZd�I���55�ԊQ��6���e��qܪ�W�O4x��AX�i�xm��F���vQ/� @j
�ć�Q�ZΓ6�spO��p�S��X�PS�<�P�#P>|G�?�1 b�1;��$!p��_�z�mW����N^���-���s�c�ev�u[�V-X�Q�J�jK���U�l����6^�z���N�d���8%ӨW�?������#���M�ɨ��9�J� �&-�����?�9�?���5��[&�:U&B0���⣨Y�1��)Z�`�B ��p���BH��o� ַ`c#gll쌝�?aC�#�6�JS5Ǝ�L�?U>�5����eQ�H�M��3�ȑXuax6��lt>ߩ&>�X��H�
Xm(ƀ(�ƈ�_Xn��f;P��G2!�d��A�uE����	��P�#A��ɠ%f��!�SA7q圏��kh�xo板au����;B��@Ӈ7��z��Kr�	Łkആ�x1�J?�B����ի�z�o������`==�Q���]��J۹�
�L:a�j�R�v[��޽Q�\M�jn@����I�әk8�H�'��"��d�b��6�<Z&�|�=�|�%��.�{wk�֙��/!p���:�VB<�ł���'��3)� 4�?_�����R? ��؉���@�Ɔ���G%_R�6;�7`߾��Z�����4�˗��ZםJ��Z �@,*%0�|h�Ӂ/K5R�m�iu>����ب	�H�Nw�l��ę�6���G�����P���gW�>�V�6�=t�J���S��r�</s�ld���Y x�Y�sg<%��.�v�۸/V � �Q��t��O"�_ Z����45p��9y��7�|��X#�s�e�u˥V��{�b�����*ik��U=���*��oo��J������׵�����r�7�H)�\���i�_�������6p���!�4���F�hB#�nr�'�جh�a�n����q��4K�-�"Sr��������8j�Ҙe3˥��]�;�w̱#����S�BUh�+����ΪY��C3BP >��je��8N�p I9V�ĮPs
AZ!��C�C�V��i��DA���y���ID*a ���E�*�F��(,������~;��k����s���������_/�!�}Ё!�F�^����?����ʃ�k�`~�����\��������f��A۵�J���͖JT�FD1�n�u��x�f͚g�]�j-�-��p��{�R�'��:�%I����)�p�7��LE�|&���[S>��(��S8|��帝��A�C�h�>��Xlbi~�z�@��V��^{Ķ��mլK�g��Jy������j%��LZ[{��}��~�)�4)V�I�'��B�Oʣ�������y~�a�TdC�Zn�y*�G �	7�+Q�l�i$����xEIp�q�M�Lo�O<t�4q<����&��$_ׄz�2�Г%#�E� �*�;��է`)�@�yF`p}��*Ĕ��0���r��B	��@l���.8|U�'������s4pﵜ[ӣ��o߶��ch�J8��Ixe�f�����M�Z�Y"�v�8U]��'�G=�{/�]ȘJ�z��T�P$T@��iGd����i�}��}�����00��(�	���&�\0	/c�jz�5e9��kG��d�h��h:m��wl�*�#F��$��g�R6{����B��J�l6��˩'ν0�������J�*��c�㈆�����w�C�1/p��7p� z�(+��8���y*#	���&�Fq�Y(Jl��⚊D�#Y��r$��g�A&6�|���0�H���r�9��W9�0�D������h��=�x��(r-j���h�{?�E�,���Y���,�oV+Y�2�Y�:,��rw��/V�\JX���L�ݪ��er9+�"���~~0j����z�S����d�˼`�[����jg4�O�O&_��f����K��f�vv���8<<��ZWW�'Zș'`�����W�� /i��AܫUy?-{��{�"�4j$$%��5��.�'��L�#3e�j�8Y%���w`���ݿO����
��^@4�v���4v� E,)��r%1�/JbGCb���K���`��wfgg��������~��eؙ!�/��s]{�Ιs��y��������4�dh:wx��܇���K��s��P����9�D���}�)��H֬\�bi�RP�UK��̯Y5V���M-�m��,;P�Z,i�x�^ۇ�<�\32���*cS�L���W��/t"4`��ɣ:�.0���
:=��9��������Z���}F��?�����2|�s %-%_{{���'�oނ��h�bkjn�b�`'QX�����>셖��Z��mJ#`�ʙ��D��~�]1�p�Q����G���?������Xv���ɘ�ke��b:�����%;|�۲y4#:=Ǽ�ϼ���/����E�PE�g}�$�h<<H A�?yF�=z���q��#f���>5/�]�	�36y�Xˤ(�V��Y�,f�B��?�.��f�B3���h���O����G��?~ꖺ�&�!�o~�o��@���������&3]rT���j����cC����Δ�o�׎>f�==~��Jf7π�?|.�?yʤ�x�?=t���f.$q�������
d�-[�£+H�bQ�z�=�ڹB*�&�v��qkۿ����7<2m=��"�H�!,��pp�*� �?8OTI�7}�fC^��}ʶkףv�s���ojL8�{נXʒ�&۹����v;q�ߒ�Fw`�@�3;������q��#N'���E��f�Q:�
N�@[I8�
���
�g���
�7=Ŀ�ᛈ�l����v�RkH�;|I��KY�T�ɓf؆�[��D�56��8�b��e�X���S��)E��:F�i��!AHTAx.o)�''>�/k�3?c�L��!������d>�
�B�f��zh�}��o�B`�ވ����G+�f͂������R{�e/{��$9�6V�y�R�d���8���9,�xZ���X��O</U��%�0d�ǆ�4.��i�z���ݹ���>dU��J��V��KZ:�b:���������[��٩�ٳ��O{J	�����U�S��M�ld���#����B��X�N��u��7aȹ�>Gg�4���RD���5�ym3���c�u�e&��S}�y�_d�
��)��i�4y��=4��t`8�u���J,@��<���=���(�¿r��J����`-#jzz�F���������>�;u*�&�yt�����G+�K:"Mq�^��^��ߴ�&
d嬘�z�*Ijjij�~!�7�_o�c�Y�q�;R�i��z7����&Fm_lJ�aB�9��C� 0�}�$�{��>��������:h��)��oHc�P,Y:�jm{=%ɋ����-��>8|�?R�/B���Ĵ��8�t�OC�ۢQ;Q�����}��Ϲa�7��S��$��F��ty���+�T�ui��5�wcV,e��u�57�؊U�,f��Oo(�G�m�稱��~��?��p�(@�ƴ'e����Om��Paޣ���D}g���%���T �����jժ-\�ȦO�i�M�J7xe�}m쓟�����Y�q�uV�>[�m�����Z�
�8aV������������y;�^{��?��J�R�FsC�]�b��^w����$�P7 T�=��s#D�j�rS㇘a�ˡ����|caRu2Z�-/|ڱJѱ���tٱcv�H��v����Z,D, ��=�e��+���T���s��
#�w`c)5D/����y�_�.~_a�}E��2Z��#�����xN��������>/�y�J+��M'�&mN-=�V��d�w�
eknj�dH�:d�!�1V���GA��د��Z��l��	����G��?�yg�r-��|[6��B~����:w����}���㌍�0�^��ټ�����Ŋ��=�ȣv��
�CB��.�?i��t�m�������xOo�ug��B�Rɸ���/�+.����Az觶{ד�L%,�ΈU���ռ�ґ�ݶh�{�^7�%J�I��ۭ�B곐�T�;������g�d|l��r�$��/@����U*v��k߷ݣH�u���{��6�CcOz�r���>Ϥ��(6>�����ƣ�Ȅ	�|N��Tq���F>/:8j	����C���b�97�g��v��\�_m�<`kW�g7���d�j�l��O�j�nt��n2��3C"��D@!��By�������
�l�r[�q��� ��@�6
UpaB&|���|�j�(��jκ�qő���sߙ�6;r䘭]���ѓ���n��K_��=��9�i_^�u���oV	�ل���}�-[z��
v�}w۬����T�:�a�R�q�%�iJ��;U�W��k��/>��� �$qू#� :,�Ph����8�}Ī)K�O5k�N򪞅b�'�466[[�A�����=A��@�ޣ�����o�z��$y1.�K'�W��;�E4u��te��2�yM�bcC�\�9{�e����h��%���=6X�9�ۜ�X��6oZm�*��kV+Vm��%6k�*+V�V.��Z����ӂ�G�� ���G�b�[�ƌku*�� �3�u!���T�_�?e?8�rΎ����`:;;,I+�xh��Y=|����g-�/����fϙg�x���;�5(���>g��m��zz�����[�O�<���G�q���������9z��zp����w[��#�y$kK��R��Z��7�<�4C�P��B��ҡ�����]��<l$6E�p��覧�l�z��b�͚�v�H������}��W,a�;�����S{��X���i��U��x�Ё�+_��]r�e~ppӺ񢋶�&�l���/�9�a��&�.=CY�r����-�0�c�S���+���˸�r.��Z~*�B�V�a-���/�t4F[y
��U����������*�Aa���>����4�Ud-���I�ɀ��i�pMeG�*(�.c>�x����E!ߌ�M~�9�����-ާ�E)K����՞Pb��
���p�O/���f�b۲e�U�}�L&,^1�>k��Y��*��b���:=s= ��Y苡�B�����2&���y[�]�W�������N$��O'?U��_�����'��&Nh�	�Z��=���Y�6Y6W��;;�RK�ɓ��v����rNM�O�3�x�VXt�G��,�}F�PՒE�?w�]�u���>�����]v�k=R���C����fX2��S������i��q�V������R�'�:��fs���OO������'�����r Y�7kH&,��Y�������;݁��4���uڽ�?d�\���Й����z���ꆍJF�a���osС�O6��m��^@G/V�OMz� ��9P��<(<T�) ��-0侀���h"m|���(�34�@ 
K5v�q+��ļh��V�ͅP�ƨ�`	�A�Q�ƭ�b͇~�<J H��Ґ?�s0^�c� ��:�� ��
�1N֌9�s\�N��t�%��4]���ֽ���u��C���D��*�%�,0"�O�흼���7sQ'���%��X��+ϳ͛WY��o���e?a��]��;y�����/��͵r������~��)g��⋼�<?
g�fCP��৒��g����}������ov�sm⤱�c�ϭR����l�v�9`k�����\���B�x�����=%S=j���Y���>���[���v��U��@�}�߰�/�`�X�����p���Y;r�U*��v�5L96:�ޮ�_�MMo>� @�����}׭��8��u UR*��%gt��J�����}����SGͪ��h0��X۳'8|��g.�����!�s�h(��h'����c��<c�={���;<�B~�֕$�ѺR�BQmz(�I��(xHs�ʀ��F#�� �� �!��Um 	"��Lt�+�O���{�nc0	��J{H *������q�"� �p��B�u��2~=�,�cM�^�F[����?�HT�%��c�\SV��������e�N8��p���u����+��P�!��6�X�p����o�8�4i>��x�ɚ�L�ISfz#u2���N�C��g7̅yt������-1�G��G�O�'���g�+�K�X��ڳ�q{��o�ʕ�l��V۽g��$��Rͪ��=���4���'\���
�U�yٮ={�'����G2Z��Po1X�{�����?�^�ɪ��>�����L}���'��[.�#]�A�G��ѡ��,"�J
�PP��8|��l43q�j���<b�o�`:~f�OX�T�LC4�x���i��費�}����&�T 5�3O�����P�\�4s���6���^�!�P9\�k�6����0c#���)o,�|G7�6�4h��@F�q�'j�*�,��QPR䖛�ޗ9lE*�vQ�d���
n����S��PU�b�    IDAT ƳH;}$@�΅��h.���q�
�|J�������o�;���X��yn�8lֆ=�ƪ����T9������2�%$������{�{G�uGC�����z�۴q��q$��|�X"�%�s��G�<�"�z�,I"g-D��kh��]]��=�Wu@��8;�[@YC�!H�f��e��٥p=����<��~������ĉ���m��KE�R��lޏ��w���2������A�����mFֽ��9��w�?�GkK����&O��η�n�S��Nul��D���T�:1`��d��/��^�җ:xP����o���'u����$�:����k�7��m�ڑ��<h����&;S��//��'�#��,�Y*�|$�D�G�9��I^ݧr�L�X�Z���9�3�|��_���_��_ٛ��&[�|���b��Ǒ��9��	~e/+�M�T4ę�( �
�J���h��p@�4K��z��4z(��c�gS�(W/*Jܺ@?��.!%zHt��*����BF 
�3o�>�����{�y�% ��2�����.�2�c�ŵ٫p�\KN%D͝Nn,��O ���Y@Q?E�ϴF<�z\h=�N�g��O�{�f�qo�N��WY<^�r)��=e�c��/k�c&��/~��*���O�;�D�P�+����i*���Y"�A��F�'��g��|,<�����8��}�~t�]6}�8ki�XGg�ˑ�PW(�~�C��ȱS���o/x���+�\j'Or���/|�N��v��|�V�YL�����&�P�xʶn��^|٥��sº�:�����8y�ʕ�%q+{S���c);~�{���&�_��5N�pҹ��ˁ���~���XhWl2{��A�_u���=Z��r6ƦM�BM��7<C$y��8j�	�$k�JIgw8�c�δ؎���;��;g�t�K��S�'1�#w�Ղ�O�UW]��� @���w���C{��"��j���E]��1����-��0�QJCܺ�n6���Ґ��^`!MYZ��q�9�w�;E��q�v���ʚ�`":F<u��$Ǯ��k���`�~Y%|�W�bQ;r���FAC�X��`3$��0c�,9��ή]�|��@�{I(���[ȱ�Ϩ7��G�,YC�LtMt]~
�7/��:�|:"��×f.O�}��_��Ų���CSC�J�|�y��Y������V/�\)ǩ�˜�7n�;~�~����zg�@߲�?�я:��<+����}h��h�����u���u�ú���l�+������	;��k:�X_o�^�����f�2v���; ��*hρ�(�݈v�I3���׿�Z�Ҿ:�ڮ�OZo�)KRʙ�o޹'i�J�j��󗬶+��!��D�s�{�8�}� ő�/��O��/��n��&w&�Y�!g�{��(�U����W�R�Y:�D2f�b�R�F+Wv�D���5wX[,f��p`f>��>h+��7�!lj����r�']�|�;��!��gy@���A�C[=r9(ꔅ	ˋM�5ѐY>��h�(�A���|>�;c D!�!�9�X�+g��|0���5U���" Y'����Su��S*Ғ�{��)J�uHj͹�"���s-�s͘��s4K5|ѳȂ���]�z���&\�R"��s��PEX���H�p]�IT����v(9o͙�>��Ng�)A��D��(E!���8�-K��J`�4E��.�8�O���~)�L��榘�C�D�O���|�i��U��(�@Ѵ�eZ\�O{�>��+���A�_��Я���(+KJ�g���I<���jլ���i���Y6G���G�Bɚ[-�/{��qc'��������;��A��3ٔf6jU�xh�H]Up��ۅm�9�j�����O~�#;��a�b�-�;ޖ/_a��l�Y�X_߀o��[�V�?8|�q�I����?���]w���x<l��f�\(���G�;�k���Y���T�fU��d��h?GtO�,��д"�$V%���U=�|F�d<�&Z?4����N>�ʳ~�S��tTϏ��\2� �Ќ �K@�"��B`��}��ph�'�y8�&�$� ,�.-|$��0�9��LBp��"hq���c�)��cf��G)cz��\�3�G �<��3���Ҁ&���V}���K^����p/��K#`"K.v�ʘ��ʕ+]��pD������sM9b�����d���5t$��{�;�\��9���5`mn|�y�����x������e�l�B���`�����݊�8|�	��˖0�Eђ���b�X�
Ţ+J�Z�&O�i˖��J~?�%�I���Wc#M[ʮ����u@�'�����W5n	tYV�=B��[�E��ﲥK���wn�n��~;~�;�)�BH�̙sl�ʵ^h2F��Z��o_��/��t��s��!0Z=6�Lu~�u��i�F����Bo�́�����k�X�&L�ds��3/�M$~,�& ��X���ȍh�lG�I�r/�o��o�q*�tp�}v=�����I�Y�R�)B��ԩ�=��V��_f��˂�l��V.#��8��WB	�fӽ�5�sڈ��9�����;�0ǯ�إ_��W�Y8�D(���@���>g�|�+�
 ӵk�:� ��CMH�A�O^UNB�+�xrσ%G����kD�5k�g��0gPvX)j�~�m�����6w��hx$��A�%�C�@C� \\��B����"��p=���q}� ��? ��e O(@+ׄ˿���z���گ9@�RB��<@�#��Bp���[n���F�+���A(�,W, ��A,� ��]����g��,��3��E���������}rMX#� ���`��=4[��ૈ�D�)�oO�2|G���[8o�-]�Ъ%:��=I���R�f3gͷ+.�;W�����)錒�X����=uʱ��y�E���u���/�gy�����\�
�8C	y�k_m��u��\(�Ѯ�v�P�𠱡�.\lc�O򂊍MM��?�/�v�ϕ�h�轢��^�4����$+��~P.��W��!�6��M�ߟ�����������?~Jq�lT6?}aqS1�
�\���_�ʠ�)� ��X`��\|z���_�O<hǺ�[KC�J���ͦ�Ix�۾}�=��G<f�B�C�jη���
����C����׿Ձ�g��׾fO<�sOhan���@q��!����t8�� _��v��)�2�4y@Q��p,�\��ܓ���'�=�y�s� ��.�`ܙ�\�w�֭x �	5B��9����T�y��b�/�uh0ƈ?��lXH 4���S L�}XX '�A���l�F�'���	��!8s�<#τpŢ �����ٯP��9����y�#�*G�o��o�}X։�@�s/�k�6�����,����1�&�N�}Ü�̿���ꂛy欈Fb��'�)����f�G��h��v4���Ϫ��m�ƕN��I_��j�wĬ�e��]�Ɋ%B&���|ɝ��7�C�;��n�[��H�?a�$Wz��ST${�3L�?���Žy�W��J�9a�Xߋ�Jy��Q(S��[=���;��g�5g=��h�6W������ji��0O��!�K���D�������^�>��x*�>��'o;w��~��v����2�i�p�ho�xh��o��MZ �D����}?�
��hh�̑���l���Б���Ү%KŃ�_���j���{~�����=�B E����B��ac��‿�s����::� P|ի^b�=�<�����h� 0g^8$r2����a����G ˈ�Vh�h��6 
��ÆF����%�!�   <րC��"Дo�sO�t@��v�o4~�eВ0P0��� P�V��r`�,��5f�h�h̀>ό���	B >�3�@�4N��5��'�)$F� ��AX"�����Cb1�>�����D�p},&����A�#�{"`���9�^��.�'����#9��� b�y&4c��Dp` h�OΎ"�$ ���;|)�P,���5K<cߪy���Z�a'�P�z���u[,�i�r��u'�' ����?�1����,�ٳ�z�7�6���|�c�R�ϣ\$@�yϿ�.ܼ��iTidM�p��v%�$Mŭ�ʺ�w&!pVW��b�����y�p�O��Or>�is�Nu�9cƌ�C���lX���~Sf�Y��ϡ��&����CE���� ���Pa��4��p�n�R�֒9oP�]���x� �}8�2��,^|�M�>���G��PB[�N���k|�2'X��O��2�(���������{ #a��|̫,$@����3�I��������Ƽ1���
���so��f
�:tȅ��ڱ�rJs]@���1���9�p#���c�q�C�kG���P"$������=� �'����~ m��S��Oh�B����F�h�PiD�(D���[).�`yp=��8q�<��ڡ�h�X8�)��E�@��B8 �/��s!�z���j��=Þ�o�`�Z@X#@x&�-
7)oӦΪG��9ڇ�ΔQ�$����R�Z��W5|l)��B��1c'�KVX2�h��R�Wt���op���|��.(YC����}���d�27��!�."���f���`��R����B��X����ΰ�E���Z<a}�Hk�^g5�_~�����j8�?�$�v�"M<�B!;�~����t�oEˤ��TZ��B��_��_��Dy��C��h�����-�q"z-�x����U=���Wky+�؞}O؉c�,ӀI�������j�,�ޤ�+$y-�3��V��h�?�q�$y�I�1 �}�� D��PCc( Q�Y/Om����������I����Y��]�Ce�2��e�?�C�p� �	x�
#�@c:s���4n@P�|O��1&��[�L�#��z ���@`��h��A	N\�ﲏ?ό Ch�>��2V���%��7�G��X�D�H��3
I�E� <PMF@]{T,4�dyvE�)Z�9�|ȷ�ȗ(��'�s�gB�����{�L�nY����O�����5��zl��e�y�*���Z�jD�4�،����ɳ����C����k�t���y�5��S�7��>*���<ɡ�{�_�A� �a>�'='ק�K�ۛ���!D���+,s�9E���r�����2���=|�]񩞞�7�nB����Oo4B:}����K[?8�нG���f�)'���q���9�8���X@1���5�{���G�R�Ǣ����s���ai	�fh��n��v��S������>ف��b�:�/�&R	����11^LN�����(h�������"��?h/4>Q��h��1�����%=��b�a��
	�o
)0E�ֈ��'�(��Xt��U�d�H�(�C�T+�� `|Ou\��>�Z��\GQR$����r=��M֤"�؛\K�+t�g��*���r�!���e�!D���h�|NJ��#d���?`�gEI��<p-��n���:��b%p�}��i����y����}�+�АIX!�m�/�u�.���_�ڤI��${*=�jP<��;�G��@�<ɋ�?
������8�U	���U���B��u���@���38���8��h>���i���@Q��4�)�&_{��f�������I�����fU̓<�0s��җP1����7eZ���wP�OA�
�xk4A8Mi8�������>��G>2�@h���*�v&��"a)KZ���L�b]'xI�b)�<���?l���'^�ڧR�;(�R��p�����p�vc����b>p�AO *  �Qx
��ϡBbJ����7�����[U�l\��aN�	3~Ɔ���@B���u|�4~w��+|
��;��X�@��*?@Bٰ��W������)M�����ݮ��{K8z_龾A_��q�����T��br�	�
G2t����N��!����G�Gs%��s�̫���{�4����SF5SM!Q�Q�$���[��8^`k�,�t�jTM�C���KmּU��W���d2�)-$t��hL{G0��sS��O����� e_�w�5�Y��`-�|� <j�� �J�=���u���zC�
�J���B)���z�s��f��m�>�����3j�5����^���
~BX.FA������]*�tS�8yN�IT�d� Lp�*(Հ���o�;~0U����UճZ���=Cq7�>5J0c2;z�ö?��� ��2����{?[�D�����/tǫk6�vc�\�y�X4�F�I|���s�� � Z<�,��CX��@ �
�s/zB�%��i�:P�'�4DJ�LS~���e�&d�E�1i_|A��4Ƭ���"��rUn�������wyN�/��Z�l��D�B��A�/E���" x�Q8���e �������J���a˜��+!-Ag���|f(x�<����tV��Z�B�������B��p���S$'g�-�իϳT�j�R�
��-\����_c�J�2���C�Fē�z��Ԩr>��W/G(Z=��,Z��!�'�H�#��u��ϧS��T=��s���)�����M'�<�s��030�'b�$n�
�w+�/�ԁ{+�U�6�{��O&��4�W��{�ő&�CqzA��E��u���ٗJƬ�����s�>q�k�P��H���G��w�o�Y��]F�9#��� �5�����s�n��R������C��� �04�Q���H?��<#��sv�P:�kp �� ��f�=_A��m�T���z)dt@��ӜųhW�\h[6�6����)U-�j�9�۬��󗢇�r���p,|����`�̠q�T�,�`�?���*��n��di5fBR�W�> i�I�=�B��C�����ʭ����y�p��B�	� n�bg����!rE�* ;!��<�B�������H&��c6 �?�hrI��a^����:���O�c�d/�J��il����=���
�PŇ����_d�f�䅹;r���ND�?��NJ]*�ϸ���,����m �_ڰ��у�\�g�5��'����/�n~6?�pc{��O�R��{�nظ�jeJ9Sч�кcl�����:ަL�a��YS�8/�\Ĳ��W�lx@������9T`�4{�9�S�Ƈ�#�NTD�<gIB9��"r�T>���Z
V�5����OX�<��?i�|��>;t.��s���?^�`�U}�tTN�`~�<��S�.y%P��K�e�e�G�;�F�Y��l�-( 'Ǐ�P�UG�v�P���u�I��Q�J՚[&؞������C=�	Vb68�PO|u�p$�!$��5�\��Q矿���0�I�����""H�h��Eل����^��p�b=Ȁ;�q�z4ƿ����* I^O�����C3�zd�mӆl�����ސ�X�HDƊ嘍i�`7]h�<�C��*UK%3�h@��$�|��A�od�K(��ɏ�)�Q���N)5�y�B('Ih!h!j$�ǕM|�жi�Џ�7p?K�$��J<���3A�NXA�w��\� ��0�j$�}���$�37�k#̐�I��Åz�����G�\���7�-V/�[�O�l��'��{�%�S�&.�g͘�tV�p�����f�����t�+��ꡉ8��w��ͳ@-��I�l���<�8;�� 9N�{�����ϥy*�?��C �vklHY6�m�V/���ά��(
"� �X��Ŋ�3Ѷ\x���!L
�'I^|	�-�s�\�5��;���9O�����ij�e��+��R*{���	-G4}�ߛ0�&�:�O�2�/����{�i��D�T��o�+�����'/� ~P���N�B�#a!� J�@��G�'`K4�����B�CT$o�    IDAT=��5f8��'Z�����UK���֫Ikk?b?r��z�I�}p�͟;��1�	�EG�F���ybŊP'��@<8B�������AU/�+��{.��sm��טkY�RZ��ϵg��2���O=,r����CU�T�,ޒ-^0Ӗ-_d��P�Y2��`
��?�2��l����b��/& V ���_��C�dE��E�I�Q��a��b�!(T%����G
������������ng�O=���n���:���$/xp�RK�)�Q��G�"qy)|���(� Z@��(���Ђ밍�Y)"M�Q/�ŦË�
��[�Zo�I/�L�(�&V�ZKZS�D��/x�z�@%[�p�͟7+d�B�h�K8y\�<�-�08^�|@�':ģ�Ik
��B�P�gb=���2fEJ�Sʌ�tT���2��8Nk�Q�9���:���Z�2��%S+�<d���P���Lc�%S���<�*U��:�� �zb� /�y��Y⥈,�a���5�.U��AqW����x(9%"���g���K0傥����O�4����G+�P����h�l�F��S�jH���-t�pnii�E�e��,�;�vR�66��uF�5��Q�o�j�x�I]���v's��}m�����>K��?Md���d�}y�1�'��Λ�%��//�k8�G\����o
܉���\����X1��p4ro����}�=���ϊ��"�c~Jy��U3�O�����>��t�Ϥ�V*g��9f-�)�2�+18�A��ĩ�f�z���cA�S�z
0τ�=�aťpVi�Hi��E�D�Jm(d�L��ǒ��CkS��\�ԦN�l���>Ι��<�4�87	���{��4N�R���U���b��v���`��fO�m��_�9�f�E���MJ��kRH������?�I�#�H�����iq��+��n�,�pm�6Q��?b��<i�l�e�^�ө�QJ�'v�c]����gΜn��~�3F�	��|.�WQp�����_q�K9���@��p��B�3�����g����w�OQi���?3�s>���:E�-=��Z���� �C5Oj����9k�]z鋽�o2I&P�p���!ڇr�p�(e仼���p�3�T�q�?����G��	�$'f��6�lkl�0���X�ʢ{���?�'�[���B�D����Io9+9��K:WC&/N�J(�If���+^�r�0n�s}D��S�N��\2�0Ƕo��}l	o��%�dh�
� ~�EI�UGvM�̹t���JV�^��b%۽�!��M�Ȃ��|�7N�f�ut���&%~��U��G (!e$�׭e�~&?E�Q|%J��Z��
@8ʔU���� ��Q2���
�hR
�>�@�E���~r�X�6�(��CNa�<��!�\���F����I�o9�d��}�C�+�\t"�a���C��d9�"HX#Y����"K�<������h�g.f�]�|*��퓴B�7�wX�ܬ��n+W,��X-�h�bŒ���[(a!�����;`�&ݟu���6Dӕ�^���W؟�ٟ�Y�B�zq~ɘ�ҭjT)L�(��m��\��Ək�=��'�0c%8�����;�)���`��fa+4t����Z����ꎢX�3M~�_do|�묥�1X�>|�v<��u>hM�F�=w��w��:e�KUK�3��J-6
�!P�v=un���S%�M�g�?��O�#�xp�>��{��ah_�x�v�z�N�8`�B֒�%c���IKc�x۳��{߃6�������i>2����hN!*~�vv�u�ɆV�3�B��E	I@ոK��(� �����åB����G�5%PD��k1&e�J�]	/�[��響�
�IX*ƛ��B�{�:�k�\OUe��7����s�R��e)Ei���sܛ�Y��ҳ�7����SB����5�	�_O��~�O��P�t*f�B�mް��o\a�b�ҙ8ͳ<ο/�9�Z[�ٺ�<ڇ��yXl,P���Tۇ�Y{���k�[�盽�P�-@(P��o��"�٦t���Y�\�\��k����<��,��#X�����^!V�>�
�P�`}O�'M�r�Y�u�֛�{z�=S���$��y\�)S�7_�*����V-Yϩ���#?�'�|�Nv���f���/�bp�]�l��^��#` �������
�S_���ԽA�!���fΞ�%��4
�C� 7R�'����	�9u�N�<l�~zc�V�X�XC�kk;����Bm�~(��}��3X��Z�lF6;σp �pg�R߈�a�J�^�q�?'�U�+����Ł�����Ɛud>)��f�9c�GF��!sH����q]擒J����z|���N�Q�D �_�� �}d���&L|�^�ʳ�ٽ�AV�E�����B�j��{��� �oX�� sĵm|Iܟ�9撹C9�w�&*/j�L�2�+�j�x�$.�mP�_�Ϟ�<�G�����S�e�r[�a�U����$�����i6a���I�@��垓!䓤O/R*�y�k��G)�����y6�d��A������#�@Nb)3�I���K����{�b��{m����s�c�굶v�&���%�Le�;��fh���BEÿ��ugga��[?���s�3|��aH� ݛ�'o|�l����kk�i?{�^���MQ�b�jI�!�j��_�%KWٺ���9����}����)�P�p��+��~͵oqI ��<hm�G���zmr�U�=�޶ݎ>�!��$2�&ۻ�34sɖ�ݤ�ϬuW����q �ď?��mkmE����u��9�S8(<֍�u@�������=���T����>�`��6�8�i��e� ~��O:�p㾔� �ɑ@s�z����cԴᙼ�s<X`���Yփ}��!�(W�㟱"����������C�s;�^MI���O>Z!�{�Y�ʝ�	z=pO�hQJ��_��"�3.������X�p�wXc�\��&h �%�����5#y��O-�b��3|�}⵼��x�fM-m���6v�T��˚�.�֡�C2c���,}~9��\������;n�Az#�����9�;��B��#���<��`A�R�q�i{�ч��'wG�1�K���z�5���V*�l` g���?��Q3�a�
��{����m���~8�w����Z�Z�7��Ͱj�h�>���������`��KK���w>W���S��_��lŮz�[h �]9�2���� ��y�k�>��O;� ro��M�D�i�=(���?Z��Uc�I&,�(Y���־o��j%�P��\��G���)�?!��_�X-�FJ��� 	��j��@?�Y^��KD��h�<� g�	 ����e��?��?�k|��?�/�@�i:z���ŢMQ�N�� ��V��F��É��`.Y�@G.�=�3`]L�:Ʌ%�)����\��hX.T'eLX>T[���vN�̯��9�K�y���?�k����;4|@��`�ױ�G��P�Mj!!d�/h@ ����{D�QdA�r�
?t"�E��BbL������g�UF�}���)�`���Z��֭_j����9#0n��l����a�Q!��]h��D�F1���:0f�����Vk<eͭ-���WzIg�?���X��a�{�ö�\>�O2Q�#��m�欄<u�{C�|��kv���,�����~�-Xx�o��|ͅ>��|RZ�(�svk���?� �i��ٟ�ɻ��a��}��ٺ˭Z�Z[�.���]��Y���v����f�tۖ���9|�2aY�K_[�G( 	��}�{���ń�۶�,@��06�\ФG�},n�Z�j�y��v�X��k{�
���
�����q����M� -6�G4?ټ<�f6���ƾ�-Fh�@�2ln9����̛@t��j)@{�'?�@e�5Lj5�ȸ/��T��µ��i<���+!r��E�s��d��C��-娱�кyV��5�y��_�6���ͅ@���u~��<��'w� �U����b>���p=,�xz#�Rv���c��+Wz�4�{
���PE�!X<(X!������e/1G졨������ь��?���D�V.[`�6,��J/x�����Y�-o�V��{�s��sJ�y=�9m'=������s~ޒ�}��wT�,`����+�	�|��{��߶���)T�N���o,�Z��}V*Ǭ�x��ʥ/�K.y��3����ӳ�i�r���=��붭���a8��DC�9m��p���J��:q�~��o��e�������ug��R�ӝ����l����6w�b�r��g��jY|�EW�q�U���e 0���"� �5����DȌ�Ex&E���:����y�
�~�E��D������i�_����
�D�'��.~_��&��w�.PD���`i^�3���IVh�h����g�xa#<�3 >��(�CA3Ѷ��];��� ���}����چ��h� ����}$˫\)�8xa�߸?��3X*_�Hx�G�((��K_�VԞ��#�lX(T<廔�� ��Iz%�	j@����}�.όe�����)8�y߳k��=#�g>��\ ���G�T�'�Wq��zU�P�'I!�ꀭ]u��߰�҉�F#��Y���u�H4[�d0�Xܳ� tѢ�&g�g~���>Ŋ͘5ӕ��v�g�Q|��P|�s��_؋�S�'��c?�x�-_��&�c;v�E%�$䥬�7k��t���v�D����`���w{%�#�N:%�s{h�?^��?��������y��m7�`�I۷�q��[_����V.�Yǁ=�M�S����Z��C��ڎ��KVx�T �k�Q���w%�GQ��b��C�븃D����>�P�3 "pJV�����Nkk{Ҋ�^knL{)j�留�}Z_��`i��l��YV�~$�a�W\?T�ҥ��8>����^��Q�]8oh4_�X>80�<��&�"(&N��3�	���C� � f��C �e_s�N��v��2� &����ϐ�?��$3��j�O�<���������G�:S��b]� о�7_��^1����h�?/�A�#��cg~^��K��_��S��茙�&X!(<B Z뭩�ѝ��
A�傰Ta����������B�Y�*���N^T�ݸn�mش�j��OTi��V��9K��������4y5\b�CE�������hwkݣ},a�}�����7��)^�q,a�S�	5��X~"�9�(��{����a�2�8q����J�Q�L�-�-��]m^|��'g=}y����ߚ[�Y.[��|�c�Ѿo���9��O/�r�Gz�{�:��_�7
Y8���Ʒ��g���v�7���������|X�j%i}�y��+���w���e���Fʣ��������B��h� #��Vv����v���@�T��/9w��y��;rp���V��Rλ6���X�ہC��{�L�LC�
Xϛ7'���k����+�ꪩ�%����'������n�Mp�j<�g����;��w�P���] ���,%4o�V�Z"�`'�1 ,C�i�p�{�X�y��o��8��>%�X#iϬ-�`�<�Ȝ�7Y�'�{X>�=����>��<3���������+��F�0G(���w�� �N��Rr��ޔ^{I���B�OE�9R�آԠr:Ȣ B(�i�U	��8�D���c�#fӽ�?�\���(���O���[�fm�ʅ�y�*K'jV,����V($��a���0�����uʜתa�]!����٩>4�P2� ~ᅛ}MX�T�jemI�"�G�����??w�z�~t�7lŊ�6}�T{��G�Z�'/h���,�h��G���d�'n�L�����ܳg��&���ׯC���_����~�<�d��Fx������w��55��Z�ٿ��?�E�-m�W����!y���~��~�ʵ�=^��.�
�L6a]8�?��X�K.��M4/�M��p-]��7����nΣQ@���Wԑ�{T�|�������U�$%��*W�6n�4{��6��COZ_o1����m��6w������r�у��P̊� j��U恟�gW��*��h�\W	[��G��F���j��\ �\��o�D%W)�_��Z����
��}�[���9�џ�R�38e�)7@m�J@SG�~݋uT8��y�3��5ŕG�A֏��T)�?��b�?p�T��	�g!c�9�H$���O�mUP�/�BC׋�c��14���H,,�:y͝��N^�5���Ջm��%��o����:M�ן�1�&��~�R���{��J=�'a1����[�p�Z�I�я~�[�2.|?(������s*kN������g��g����1}�577Z{�^��(��T�1{�g;-�i��ǻmݺ�쥿��Ǝ�d�v����S�N�?���[g/��F�`�1aM��r�6[�v��,���ʀuu:���]����J7ہ���y脝8U�����\�����)�8����H���щ���ܻ��ݩ*f�/��hn�t���Ås�}�N�Q��s�
�>76���L|�����x؎�pb��Ϝ19�i�*pÃ?�*�#�s���f-j`E3�=Z�Rq *��<)��M���P�: #Z/��?@(�s}����=s����氢a�!�=�/�&��X
<#���+ˁ{�ys}�+��s�;�Sy�ų�󀇚�3V�����%$��3�¼���{pO�Y;w˴�V�,��ʭ���7��2��J�����ESro������i�E�:�Z�(���~	����?w�i��U<�w��́���W,؆u���-k���'E���%l�l���j�/Xn�\Ś[�?�Y�����[��Af���!jg�	��Z��BAOr�yvĬ7c���p��+���'-��B1�:�3ꊱ�-�c��?o?��Þ�՛�����S��w�|F����l@��Q�&O��K�����N�b�8�P<ekW���\s�UJ9+���c�#��Ȟ�ŇO��	ո�eK�(���.X������㧲K�����+�� �N��p��׹�@4�����pM����f6���-�g�'��b�ϓ�0)S�9�{o�=�}��lt��l���6s�3JZ�� ��p�0Y�d�8q�/���9p�lv�`����������9<�CB� �t��	��3C����4Y�(������*x2��a�������<BN<�����rc\|�5b�rƁPC�#�/������@ �(�7~|!̓'dM��kϸ���S��d�TB�H�W�>�a~� "�D@/��f�j�0�`��٫Ap�7et�������b��,C	,��>�KSԂ��W�N��ГV++Hc~
��4�o��L��^[�`�-[���P�������y���<j�B��O�����ʁ��k���k�Tj;g��r�-!(�=�S�e��Q��3�l��U�}�־�������',CK�B?��ez��6o���n�fkjn�����˭_�g��%dߟ�Uo�r����+>������8O�f�KUZj�<���T�����~��ֶw�e�h	w�,�`��۰��;���,.�@4HT{��%��F� ��c��M�1݋E�� ��!���>�i؃A5���=�i�|����!b�b�s�X���V,�(ڢ��'���5�>h�42�q��
-��w�r�g(0E���n����K4Q4~g���l�� a�1�e�XHD�`#�=959��4s��7�a0�����D�0��:"��y;D��	��B���p����0v7B�8k��e�#܈���K4 �{�
 �m���5'��H/�V���A� ��׮Q!5��8h��J��u�Þ�E�;�'_�T��@;���ח��U��5foHj�D���	0G�}$��\��=b    IDATG�ߟ1mz��{���������T�p���^��S�*�����z�2��6~�Tki�h�}Yo�B�x�O����H�T��Q�z��#��"�e@ԗ(4YF(6��Z�`Ǐ�����ܹ�:vX:�r��YҦO�iny�-Z��b�����/~�KFU"�Fz���?ra7B�b�@��@s������:�?g�d{h�`'O��G:�6q�T�>m���0�
� �qڢՉ{�@�9d ����w~�@�8��� p�1�f��gpͬ}�>{�G�����U�9�N��Œ�u"g���x��*U"�ʶh��={�����5���c�U��o��Vki��I���p��Y �Z᪀. �Q�A��{r��	r� ��L��;L�� �ѦBݓfP"bEEf1���y��Qr��/͔�� >�q�L|r-7���C# ̱$�=������N4"< |�|��)��%�M��~��pX�V���yf��1��x��rҨ����s�8\W&�0峚	)-eq�Q�_�蜨�XV��Y~}G�CV\0�0	Y.<{��s�����P��7�v<Q���36ab�ūeKg���L�<O�P*ٔi���/���4��>�XҊ����T"��n�5��jj����'c�p�����|D��(�2��o�iӧXKK�u�:aǎ���9y��Ek���lμ��L|���;v�W��ekko�Ʀ��p����+F,�������F�m��������
[�t���9-^E����꤀S��O#Z�*5ʉ���&�Xt�.g`А(���녺�.p y��H��fO>��>��V�D�f2�Gi"���\���{к{�Pn�g�3g�͙=}��	��4���Bp�]]�|��PG�k�dx�MJ�����? bM �p��������NT��ׅ���a�p1.���4l~b����.f6�:V �6��pFx`�Y�ϸ� �p����j��u$�@���s*�-���`a<<'�\�
Q_�����-%�ː=��QA8��9a��o9��KQ�;�ы�����×����t~2�*�w&�"�)?�׿�w��`���'F�[J���p ���,
�u�{3f̪w�:s=��\�ٚU�m�U�<x��$Z��^7a�]��_�^M�c��A��),2�����@_���;�|=�?�>�x�;˺D��x֐u�|�+��+�!(����l��M[[�z�Fj��FX�߼�۱�I����G�p���)��;+�}Fn悃,t��@�ĭ��j�9k�4��.��6n\ocƵ���d/c��'�w�s�k�Q�5�Iy��k��B:|0�OM��W��8sB=���u}��V��;~f'�z;G��	�DXa2����~���!��@ uP��ϡ�H�l^�3P&���}�k_qpE�E��	��xf��d0��M����{�s���3��X U ��2P$� n~"��_���9��\��.L�Do0� >Z5c"��sPX ��'z�g����7�@p���\!w�5�8�@�E�>'���Rh����>� �b`��;�[�M�	��H/�.�0@��v�sF�xi�cBԌ�'��Ⱥ�x�τP�rGi��>e,������ʘk���sO���@��B���I{e(D�?�$�,
B�4iJ��^�?�N��n��ev�5���Z*�L"c�r��u]�w6v��Z��� F!�Y:�`U��jN�p^?����A��NJFdh��V2�{��nͣ,){P��]�K�㖑Q��]I?X1w~�N;x�@(��sX��b���j�Z�2i�gea���8R�#����K�ZM��%�Ny	 b�d?y�7���{,]o����,8��& ���������h��f`S����7Ra7�:�&>}�����FS���������?��T�
�!�J:��q�9G+��a'�u��� �E��3*MV5  ��\xm �a�E����y�&��� ���=�@�= D�����YE�p-�V��=s��m�{@�0���	���,kD�Q2�@�]����@P��C �yc�h�(? !��"���hrMb��h�0i�\��M"�9�惤D%�y< s�P&"�u�>\ۭ�tz����9o��~/�c����S�eNX�B�����J��ҳ�I � Z�5�%��q�?�f.���[�������X������R5�i+T����-8υ���i�BD�"�����7�)��66X���^����U��^�0?��^��b��;��Y�g��:8�<�´������Dw��U�EK%C2�sWü��[�ʒ����C<�)�t}ʋ��J)$	ł��� ��kj�;:,J:�	p���x�l���z�'k�U�������$�z̳�?��R��d����;R� ��4s�8
�s�eL�P���b�n�*iH�N �h��zդgNWϼ�.�Xڧ�4F��84�����gĽ2~Ơh �3�7��6�h�pW��r�	+��9S�-�仌��Sa��}$�枊����O8a,H����9�F)���h?��C�� �&;���yQq!���^e}��e���~��{�}�s/|-�e�K��B`" �h7o?�:%X��	+,�#�	�G`�Z`/Θ>�����!bi(��鞵5+��u�\9Jz�k"��է��isl���ij���B�l�J���S�롞��>p��Y���&R)+�r�V�/��5V������"��(b�>7D#y�!�h�4��M��j}\X�����b�����}����
fR�%;���j{��zCo���A
>��,H����^r�Ձ֏���D��P�#��'�[>4OBBh�7O�<�����{n��y��r�R�c���p��u�k���g�?��q��(ِ��IA���<��m��1f7��|q�q�r^lz�I�աW��(��p99��:5�L9�&����j��:�-�V��Ys>/�Ut
ϫ{i��$%����D"m�46�����N}nDo(�����XO��G�W���}�;4Hi�DXae<���^��1 HZXS�?�+�Nܓy��}�53��דlV ����ʇ`]��_���,�:8ЙX}�M��O�0Ux(�+����^�2�X�X�Z(�i�C�W�����ﭽ��~���v�4ѨkV)V��e�-Y��2c=��.^iώ�z
����	sa���ߛ��S��\�W�d͘/�rg:���9��N���+8X ^&\��H4�Z�{^<h>�P���(�;��=�L�� u͟�^�����Hl0�������F�_�%^��A��g8DD�l��B��Y" ������ 	������w���Y��S�*a��G��͜5���B�؀����w� /LH�=���V4:>�Ӕ�D�h�p�p4H9���B��h)�(� 0��VH"��eP&h�P9�Q�T��{P2h�h�P��JEà���g���c� Uċ(\?��c��l8kq�)����$��1C��S���U/��% �B@�F�Eĥ�S_��9�/�{(�ZV�@_�������#掝�����_[*�v|��I��E/r��ń��9��<?Bp0��r(i��ի9�%��4�	Ʌ�S�5�2��$�h0�/�!�G�k!�
-���Â?�/��Y.{�6mZn7� _��&�*��]a��-�l�l���Rҙ��U"D�Q�Y�����ł��
)4n�+�����S�J~]��{�H[]���[ �
_E�Rb����>�����3k��^v?��CæB�?U�L:���o�����$V]�ߞ���۝�� &�qSۣ��{��1���y
��Ъ�{�d�VJ�`:�����'�!�\
�Ā>�ihy2>��������"�	�c���w�#4X��8�8`|0g 	�K2���g�Q:T�D��!L��Ǣ"j&Q7X]|W���h� �N�(�%�b�B���1_�7@d�h��;�	�?�G\�U�q){��8]��'m�>J$����hd�?���_�h�]����O*�27�?J/�$��o��{q��g�x�R��pt{�{�A��G2�`f.��TL?���Ǉ�~�~.��%N^Ԣ�!/���b.�k(I���6uZ��sZ�W�o��C���/jum��/���J�d�r���/�CQ�������k�p����`�>)/�m��� {�hG�Z(��K�'�Gđ�9$1h�`�����?�_q����t��ax�B�Y��/
8/S�τ$�@w�0(��
�BY4`�)�C�Aw��������А��0�5F���@"̀��y܎�g�r�A�fko��K��J:W-4s��l4�_�9��V}�e��1���o�fO�����I�*��.��E2�J@��U�	`��4����@  ���P�8 �d Ѐ�*��|�*Aa5����c�!��.�
����3s-��  
�@�po��8H8�X/�<'U������/�3�����%? �$�ƺ#���!�g]�2UrӾ������lf�q
������Z.�����!�%��ĺ!�A+A%`�ܱ�]�/���|=��L����^w�y�3��ZN��
�cF0c�!DP0X;	��t����N���ok�.q�'Uݮ*��
��ҍ�_�zMj�s���רµ�C�p�cu��c%Z(�U��:�pܑ�߱�V��7f	�r��C�Qh(Q�N&�5pf�0Bԋ�&O��t�nݶ���==�?#�ӭǝ�1��s���>8xc!
Ӌ`�D�������%�@��()�;� ��h<����9|)���1^���v��n;y�Ò�rp�Vj�H5Y[�Q�羇O�%��?}����f�h�`0�n�r�cf^���ޅ  �s -<?`Kr?q ��7MH�͠�-��`B� ����E�>?4��5 }�w��� �.s!�8�l���z�j   �3r����h�|������R ��x&ƅ3ap	 �e H?����H��b P�)!�b2>r>��u����c8w����A���Љ��n!q}�A�s(�J��Y��,XM>������M����S�3{��W��khl�<ւ����{���G�����SXŬ#g��V��8�6p'�+��Wm�t"n�j�V�Z�߄�-��Y�Hᴄ5��n���Vs���Eע`����{0;��\{�gF���r�d[�l�$?��9�Bs�$�%�	qbSB���P\���$!�⊻-K��fT�h$M߳�>���=�myfd$�����5�=_���y�zֳ���փ���V�T�-TCX���gT�O��H �;FX���k��]r�O-�/"6 ���Q=����ܲ��==ݿ=2�G:��+�y�j���@�x$��[�lSo��2�'+�>�>��8m�U���ΟI0j�7V�C�vX{�~��=f��R*V),�Գ���n���������o�h1��gW��@ �D���-�' �{>t���j�i&�B��` �X�o�� ���%`�#��^2� �=��my6� ��� e (�}��z��K�P  ǳ�;W ���� ذL�2ѯciC}@��?1�U�eL� 	m�c�i�6�jG*.Yi���:�����^oL�PY�˟g�j�Pb��.�ω�	�b��b���al�� zyg,*�w������챋6m�׿�j_t�&j4�+��Ip�X�;�U�s��Ρ5��zO�w�����b�}y�x]��9��G4��iy��3��ʝ�Z֊�-\��.^�ROh�z�c�< ��w�>��	1�x�p`~�+��@��lO W�cx�����%@����޳����0'��6}�uw�z��O����G]S����+7o�FOo�F,d^��C���A��� �Z�c!1f�R�Z&I��t�^�SBQJ}���A"��5X ,e�q�'�`��g���^��XC�E*��G�7��]?��r��54R
~v��uf�
`F��k��ď>��SX� )�\�pŽ1��$��X�����R�@W���X�⻙����o �����Yx�G�`����c����B8�TAE<--tx,&PB����|���|��=��k��N:�X�B'�����bժt�(=��(2�O~	%��p�\�!��}��]�Prܧ,�����m�\ v����x2�#o��1�Yp��x�|�G��:V1��vIlǥ����546:��x���L��њc��1�v�{��Xg�#��! E�ܹ�O��}��O)f#��_�ފ�~�t:k�r��_J6n�$��%�Y�P���x���\�Q��$fG�/������|�j�:v�0j&�l�H��w��H-;�~Ľ��/`M�'#�y�hL����4�O	V����O`T�g��C�\(\�B!��{�sN�v�MwW,M�5��bV.Pf��_���f�^>/+¥m(��J�*H'~�c`�B[ <E/&wb�v�c((D��'�T��6s��`����G���~�|�q�>Fk"\I�y�Y���>:�x�G��������P��{Խ���s�9@u�X�܋��`�K������<;�����m$���`���^������ه�� &��]��K����]`aSo ��V����X�ܧ�`5����R}�����|�uJɽH�X|����"��y<�2�B��NUD��2:(+!�G&�;�
���/�Z���b��Y�y�P~|�u ̞��N�9�'xx%ހ��g�������ؑa͢������~g�w�9��g�s^΅7�K�ϙ�	�ּr�	ڧųy-V���,��kVZ"R�����K����[��l��(�� ��k�A2�����Ywoh�ٟ�YC*���?�Y����ƻ�~��+X�q��T�b����p9���?��;��1���>�Bry���UJ�S����ӯ���ۿq�Y���>f>��������I��Ix����CB
3�$��E��
�(Z�e�B���=�����h�W���p�'Mg�Jɚ���)cbx�-���v��[gW�����q�6f͜�Kny����Ț�Z�p]!X���y2���r?�G� �~��@�y"���z��"��ZM�	�D$�H�TJ4��$��p�s��¦������R�<�)�NV>����<₹GY{R�pn%�q/Ҷ�K��O%��̉�p���xMx)xP��TO���[��?��g��X��t�L�����c��b}:��#q�Jc�w}��>|/�������,�Jy5U�Z����� ����dB�(�J�8xW���+?���*��s�8~����=�W���6yJ��k�>��@\�x}���{m _�δP�d�¼L�k#�u����.������7_�ޗޫ�5׍���Ҽ����Պ��q��/���C"#�9*5�ϱ25�*~̐�w"?`���c��vr1eAk�c��p��sw=�t2�I�:���e"���y���
*k���$9�8MMf�����V���aY���:X̎v���V+��Y�Z�bs��O0y܄�6P(Z#�,zXT��/�ksg��C��h��`�t�LƯ�������
P��1 ���Ƶ�>���'H�*�zЕ�㗼)q٢K4Yd-�2Q� xn���6r���i��z�N�,�kl�V�����{l+jMV��1����_sl�A��������D�������Ρ�J\ �
�'����*��#N�	����,f���pn-bl/���#!�/�E�k�Vc;t�X��˟�2�C�"���7׌5;�F<K��<*�w$�oȦ-_豄ap�,����2����%2Y�4�;����N�����U+�iCRk��ݻ���@��\�x�I    IDATt�E��>��Ϻ�#��K��]=�%.�-�m��ܠQ�o���E_�~P���m�q0���ij�X$�6�yG�Dj�k�{�m�Y���}"0�e�9h��e˫��=�iC�,/�� ����yйm�|� ���-�1x .Y��r�ha�� ���@�i�X����n--��ˤ=��#.Q��g�Z����{i2�I�d���ϛm"Ji$��m���+� ��T)�p<Y��U!�wՕ��U�&�����_]� �_�qh����\T���������-eYr�L��D5Z��S�|��k�z�K+s/J���U���[�eK֠�x- <S��v�8�<C DupD;r-��� d@��>X������N��I8�Ȇ�������u�ߺ�)���ϖ�П���w�x�AV���<h3f�t�b-��L-Z\;�t�p��"������}�!�����G�8O�:#J��,��v�U=�.�i+V,0�-���܍��GgL�n���ם�)�B��x���/�r���h����-�_�ީ�o��g�3�����_≃��/hl8��lC:�S��J��?z����$>��9�*������?�Ο`�T�o �믻��]�B��\���bu�o�ץvP��;d�q�A�z��]�jչN��8TO�>��q��yˮY��Cf�iY�X������c�w?�%����)ƶ��_J.D�aGfB*8�X�ҭ;���{����e�>D��,]�O&e-^�ʗ�{�uC UqY�ҀkR`�����5�-��N �`. �w�EO�k$�C�9��L.��J�d�s<b$��4��c��*�>x����y(%���Ȋ��X����5h�g�q�d�s\���E��hav�2R��χ*��Q򉡼�
��=���r���=���s�<�V�ȸN&��HB��3����1u�+��s���i�?�i�S�Ѕ��r��p�5�x.	���)�0<��S�k���Vڅ�s��{�� �$V�Ž�������K�a�W�������@<�"���&��1�������[�t�0����cbC����pA����d���t���93��<���E�u�ڈqv׏dw��c���b2u�4��?��$y�V�b���NϘ6�9t&���|�2���O����x89
�o-Ł���y�L�@��Ǫ"�&:���@B��A���B�`;w�ԺzY�B����>�����ms���^�9�o�J��}O��W,d��:�Fp�[Z��D:��2�wJ2 �h�YXP��FÄF�$���Ft饗xP���}��>� n0�8X$ @*Or,�E�)E���J�.��a2�h��"�Ċ�o�&19�2��*��;�����-�<=p������Ce�M��Y9/|0E�xތ��	 �x�я�t5Ǉ.Q|����F &c�w�@8cL���`�h��x�=��� �\Ƕ���R�s�����B��9��do ˟�� 7Ή��kg_��k"������c�?��յ"ϲ~���=�l�?b�;рıh�T_ۇX��z�{m��e��5���v�o��J5n�R�Ə�l6n�r%�u~��{�0�w�g`���_��7���j�f�t�����"��2��x�4|g?1��1����@��qD:s���y��<[�>�e2$�%����=_��sx�!X>f��N���@�	N�>���o��V�<�]�|�߶m�x�>;���z��2$-�M�.����3s�"SU|6���4�L8L\H2 ���f�Q�< �Ԯ^�[��b�wv�ֶ�V��F�5_�5��%�wo�=��v��F��h���7o�!۱�h��y���C\�	�\'���@� 90�lQ��< ���H��&�{��# �dâ�\,,,"�+��)��YЋcb9�|Ѣ�3�X�XX)�`Cͱ� �(^H b�}�+Ã�<o
�2Ӹ~����ɽ��&.��<�7����ޟ㑸�+ә�)S ೨�����=� �����G��F���2�E3��L���ճc�O��O�y>��V ���?���?���YE�?��sƻ�9S��g�"I5 �3�(����wd� ���q����T<ԓ��k���˸`Fyĵ����YWح�����X�V����;$�H�$%�B�����l��ɶp�
Kgm0_v#�󧼇u���4��9d/O�1������w�B�\�2.	N���sc�+��{���x�믶���pgg{�=�����S[���7j����k���um��3�Z�y�����{DQ����=}u�[F��|�)�b�6n<�^�ZR�y�kn�k=|���U����)���Ҩ;oG���ŗ\��\}���I��Z�b�P���L�s�� �﬉	0a%���j�hR��ԋU,?pܞ����
��Ɇ�Ka��UϿb�X�-�P��U�f�(�P��)H��|Os��

���ʱԙ�ߋ�@����ŁkYu�yVX�,�,xz������aq� K��,(���� ��U�p�u�Pٖ�3�Ylx)�6,8�EZ��]�=ۯ
	���\�!����,"\ 1�����0tV4�b��d	�+d�+נ��|�'��C]���b
Xq� sWO�{9�a�0f9.ϗ�Xt� �� c��v|xWlG�>j�o�y�8�Œ�(�8k.Ԃ%p�ߙW�'ȳH�����1�����_��������v�R۰�����K��l��6}�|�0~���|C�8/��s�_԰�+���}��N����*6y��B�x~����R���7�)��*��n��6��?j��6n|���Z��>5{�寰Y3�z����vo'�{S<��8�7����nX�����k^s���a�%beoܞ�Ĭ����=�2J�R
���{��y��b®������L,'��QCrԣ�k_�]@-�D �Ky��'�?n�Z��F&`��e��n���\*����=d�����w0wsm���,(�H��������d�2��` hi���bun�`u�`�tx�,�,?��9�� �����>@V�,,HJG�i`U1��o��(րE�D0��(�@k��%p?瞻�3}ѕ�;�Z���k`q���Y�w}V�g�ǀ��҅��?���y�O�p�Tw�= ��
� �Kޢ���G��R*	L�N�g$�'�<��}d]C�K��s���ȣ�X�޹>���'�%ZJq����}�x(|`����y�#.�{Q@�,�������3�k#�>��_���y���J��n՘M�:�V�y�������c晐��F!�9i�|Ǽ��_}��LG��l�Θ�)p/�:�Zq<��^���&����֪��m�Σ���v�Z;�d���Eڑ�.+C2��|�M�8�b�?����n��.=WŉN��>�7s!����N9���=�o�tܲ��v��mͪ������u;ׇ
������:�TN���.���_�T8@�)`	������2�\l,?TG�v�$��W� �Wy��
�Ճ�J�j�׬��նm}�ʕ�gf���}�?��J����"/��?�#����\3Vu6��4�@������p\,y����m��� :�29��������"l <�?�����e�1�U�sJX� @̢�����n�kp��_q����{-N�3�[���11���\/ �W�g�f%� �b��xlâ(�7V?�f��9.�ͳe��&2��3U��.�lx7�[ �Y����<S��8d9��c9��J��$�,2�I-��s�/�c�O%τg�"ʹ�r@�f�xx�.��=��5��X$��)��:��Q���@
,�ݜ����;Pw���\�qKe�֬Yj/8�b������N�l���h�:+�Vȗ���?���{Tq4zG�I�P�ǎw�_�t��� �����^�;�`Jf��k�^�f�C��'�s��J���wYC֬�1c��^�� �:�I۵��i;x�î��[v��K,�����[n��C��zE`=tZ����C��>Κ1����m�R�;c����.�� Q�:��A����~;x��
Ť=^��3�z�D& /k_*^
r9^:�@%K +x��+\Ѡ@�`�:`r�^Փ��[��X��a{wo�d*XU�.����'�)���ޖrΜ�/��~��w�&^�g���w�4LN�^Ԅ�f�� � 7 �}�Sn�����-]�@��W2S�K9�&�hY�R�̤��z?��z�����-����{��e��j{ (1N��Иj��9�ԓ�e;%[j�^χ�=�
���?��8���zO����;������ ���H;B����kd_�)T(q � �Y�J��}���x��w�޾�6]|��Gx'�>X<�b�|����g5����jW4u;�x{Jv`1�	P&��P���%s��;)�����Jm�V�^b�?�;y�����'m���6k�Y�m�b�A�Ū'|�H���Z����j�x�c7�ڇ�>u�L����s��0�0Jx&�R��ϒD�K:l����lŊy6u�$�����BE�*I�q����=��6�i�����u����.>p�e��[ Nk�߼e�{z�Ӏ�1d=ׂ�ꬕ+�k�bM�������wϝ�i]�r�==]��SM�u��:b�r�����.r��������I�t�r*2��v�%�A��h��i"^�R��v�x̺��z	
� Z����t6z�Vk�h�"�3w�s��:��_)� ���I�A�,T~�"����lϳ�X!�: ��.e@*�\���\+�	@5����� �&%?9�~��nط~A�5�'p�3Wb��Zt�VO���X�ܯ��h��4.��K�(J�d�k�X
 �3���g�������pmx-����XR���Y�Q9�!��>ʑP�-4���1c��9'@�5J��R@����� 8cZ���?~�����&��H��Ϙ,
����h���N^��_��=p�,��VZ2�j_�z<&N�yα	�g: �C.	��D��D�% �?�2	�֗��dhlø#���Ž��c�|b���!����c�����b^��ҙ��ݷ��w�_*F�J���iu�����U��� %�@�홝;�ٌd�������_���~$�'��@]�t���~�*�A��;f���U���-�(��C�^��C��y���Z�Z���g����6zEJ&�� "V�^:?���I�$���䤙|���0A�(�������jǏ���������K��V�V2�4��t$�t�Yͻ�-��_��{*��k�v�zB�Aq���J��W� ��7�&)��ǩ�(IJܴ&���kW�W�e(p�'V1ϟg+�M��.���7ā�� �R�7�=��^ �u ���s~�'���iw}����u���&�/%�AaQ�=q��C��/���
���g�;��' U�`�B�Op�hX\�<���Pw,4,.3����q-HCG��Y���P2caN��;���KGa{��?���\7�� ��{�_�����i��Ӟ�5`��.�u�V���Z0�bi7q�e'Z63��.\l�Dƻy�H��:�hL��;��En��a����~���Q��������;O�4����-����]v׿��F&����{�b��Z�P���n���$;�v��{�?�J$�r@/�ݿo��3#����~�-'��t��9:�G2���'؟��y-�L&fw��5[��L����4�Vн�VM[_o�Z[�Y_�:��v���}5g��+c!��y�v���p�X����#L�%˖�%Ǥ����'���k��y�+���[��m��K�,c��7j�qaSm��N���G��)� �Zd���hI^Rp=^_<�:�Q�A�l .�τUr��tU?���J}kC�� 3�����A0y�K �v��n���@&zH�E.�ߎ��f{BD��[y&m�L���ST	���y�,�sX d��3����8�8}QW�^-,</>���#cDIO�PP�= ��P=�G�t�{#hK��uk�V�<<��<c/}��\����ze��3�ga�������o�UW��v ��?ng�\��@_�_������PG���3�S�$ׅ���_F�F����?j�dS1/�p����a��V)S�'��3$<��Kem\�D�p�ž ���&"����X�c4��'<N��/�ߺ��.@`� �g<d�~%��%:`�C�}�uw���i�N��q	g�}��/=a[��D�юu�lٲ���o|�Wm?��ϲ�H�s�� <�
�}N[��rOo�5#Y���2Y������k�s���-�(Y>�c�����e���LZ{�1k9�a���]�~�Ox&�*�r� �,� V��) ų���z�5��f"�J�+`�`%ԫ}F��#͖��,�1��u��ke�;����;N��e��/=|�J��fd�g��A�@8��]���� `���}q,I�ا�W��z�XT�J7��?E��L$a���(��}�p���H��[uQ�e-(|�8�hyql�~,`��⟵���!�h��`�����t�1��la�S��\��L��3Bm�3c�I1r�w<L�	),V+�`qs�LxD��.q�ߑ�@����}<+%)�W"�}��@��(����9�#��|���'�u�E��	�s�:?Q\1WD�`(��G�?���p��IXn��6n<�.8��}.�z&�]��U�)ˤ�s�Eό�{�^껇�����n�����qp�����]>G%&��ȳ��"�Q���=r��j%o�>m���HV����/b�4%-kv�h�5h��#���׽��]�֟ŝw��^�H�^������vǭw|����O��F������s�J{ӛ�h�j�*ł5��}{wz5O:��=�#��r�j=}�6}�"������PP�0�Eo����pR��A��2q�wדg��T\B$�N�T����	���
Sg春�p�Tm+�O&	�M�&[��#�u�;ޝ�Z?��f۲���*.$����җ�4��s/Ǿ��<���Tő��JR\���x,I,�ƢW�5��Q������U�< �X�Pyj�V��%/�-���5�/����i.spc,�47��.�l�_5� @Q5���m��F=D�`�J�����򈤢��&�a�g������έ��/����L��e��\���[s�7;�Y:��{��)��Z>_��	�-��X��={f�{�Y����<��cV�e0���e/}�{4ܣbP,N�w�������� 7�Z)X��xd�7EJ��
0x�i��K���k�T�]v�+���,���v�w=&�4~¨/�����?r'/+�X(���dMM��7�ٖ-[�u�a\�~j�g�>x��ʅA�t�B[�f�-;k�uu��D�7+�8I��ݨ�8���bB�
���:�k��+�í�:��y+7e���C��eqf�@Y@��i���5�B�xͥq����Ŋ:�c����_�Q Ɓ�J�~�,}��Jn+M��U}(Qr�)�p����+�l o��@ � B����j��n��nbN@�a�@7�v�;�AX�쫚F�2�M&�
}���L�;�ʊ����y*���o4�w�'��b1gMM	ה�� �{2���Ǜ9e�91h�Z�-j�`�s���Q��8S��jN�U����_��1<}�J��ŋ�Y�R���G�g�v��<J�'����Xn��]`��&o���Νv�Wi�EU��˿蜧5�o޲��{z^?���A���6A�3��3,��Oˁ����a�r��Qyoά�6k�\+US�8n�[Gdh�ؖ�@���ѷ�V  9'.9|,�����p��s�d+�7���ܼ���v��ak���L�EI�1c��+�c�e]�F!������ٳ�����\�,�_h���A���׌Sh@�PG0� l� �
Œ�Øb�3�P����L�|���Ǌ���)!��Ʊ��}�    IDATd��3( ��İ��U<�le<���ù�sa��	��"�˜!&�, �$u�D�wά���'(�V��8�}K&ʖL�l07�q�b��U�����d�r��ͯ�T��K(P��A8j��"������e����K�͛�h.�u���dA�3���빱p2�7����	�m��&��hs�Tow���y��p�*X �v�-c���_[{�W
�Li�<�Nk�r˕�����G��w�R��8m���nx�M�2q��T:�rp��8�b�W�����\+_�=q���FH~�}�IU>���KC�OQ����/�=��ּo��ckjL�@H)GFa�={ۮ����������,���&U����_�q�}d�364���+ �$hȮ`3c��R9 '���n�ɍ�N5�H������C����!@����>�+�CX��`�X�ϖ)ٹc���5�qCG�m)���I1?�@)fS�aQ]R�)����Ϝc�z����n��B�l���v��K�j�ު�bE =��gΘo���׽�s,Ny��d= �M�
�>G�����R�7_�V{٥���"o�k�:QAAeW�9�]_�}Ӧ��W��M�8ޚ��=������;�=��*�g���]{��-u���V��
ӧN{�i��9�埈k�I�Ʉ���7a�xzQ ŭ��D1Şsv׏�vK�~�,�X����[IxA�̠Ɗ���2�ؼp�1b��8J=�������ÛTSԍ��Ɔ�[X(V����~�����4�F�������w�������w4�7�lKD��ĪG#KRk�)����θ����PQ&v>jdþ,���>�O���� ���9�Z��k�W�q��^T�T�q��it�*����?�w�aI��
A�#`��QI�[�ϭ�Op7?�kk�[a�6��Ze�j�UJ9$<V��l��i�f���ן��x<.J>S��8�;��٧����3����߱��\ڍ����9F!:h6���ޕ��w������gKsY�	�%�Ugj�������:ފ2�k:ʍ��QhdS"�ͩ��
Or���x�R_�\�[xJ�����U���^�X�r5>�w��f����/�8~�%Q��!����~ ������]��Ԑ�d����Z�&O�a�w�;|���2^�%Ȃ��NYc���Ͽܽђ>@A� �C)�\X��we3��A��Po��Fߗ��#� f�U�o�Cy�Mݤ'�x������Ko�tz�H����]��M�<GEtǠ�%	I��E��C�t�2�z{{���O�
�# [Dȣ1�؎E�Le��� z5s)נG�����e�ןe]x��}������U�I+�)�7��n��-��>b��������K6��9-����ɖ-Y�^W�ҌA�*����爸$��y���z����&M��m���m���~�۾��t����à���{�0u���{�m_;y��:�o����a$ڇ��In�/���χ��^ld��ł�=n|hP�T��g���g�a�A��EF�/^8ٗL&0A3,;t�X|(%+�a8�?�붣GZWW��u
�T������.����>cV,T��3�r��NA�i��>�\�G���� ��3�c��&"��J�%H�$ aٓ�Ż���[(E�( zz����F���L#C���F���#m���,]�؟8���N����u���f��Xx�7d�/@!�9�^��zw�(ܛ��p���}�h�o���]�ܥ�I�?m˥�%��mʴ�6q�6u�l�x�Ű��U$�<W��p���_�B腲m�t�]w�[\�D�B�c��k����T]&)��d�޸=HxQ��B��,޾�^����8NC6����YG����X�V�O�>��;n���s>�=��ӨŇ�������+��O |�{h���Ui��cM�	�y�*�'����PJo{��<Y�	"����8zsg���K.۳w�l�ci��5ҵ+f�-�v���@�!��4v\R��5*�h�_,<�r��{V� �]C4���
P5R�0�@�` ���ᝳ?��{d�����V6��ˌ���Q�A�@]Я�r~���&su���A���m����!����9�z�=�}Y����#*U�^ݓ��|�袋�f.Á���s�]bm\�%�)�H�V:3�.>צ͜�u�JU�� �Hy"�'yEy,T�$�듟��Z���0���?�C�Kt��xv�R�@��˳�=`4��;������a1�ܳʐC�])�ĩa2\v�� ����Sq�/h�8��Fo�`�EE�"-���x�dM2y���O�#� ��=Ǻ��Ο	�d���YC*i�b�R�=vؚ�m��`�/T��7�������T,A�o-�nՓ�<��>�k��Ac�?i#�O�7��L����"D% �ÄfxY t�P<:�<	�m۷{�0�' ��l��>ۏ�}��ӄĵ��2����#���k�������V�^�F���G�g�>x&j��v2���`�?��J����͘�6��[��x�b���[��9w��SU/���x�Y�h�Z˗0�2f���d
'���)�h�nN�,��������k|��dqkjhp��8��uq�м,�F.�� 	��àO,h��GH<�>p�ӦO�����O���WC��?XQ-���>'�?�(E��cM��S�f@��M�H&��Vw&21QV0iFj�k)�,�IXS6fmͶw�V���9H`iii����r���' �MM������g�M�集
�R�@���ˇ�i�9��rI�b%3��� Q5O7�zD��*�xa�3V��?��%xw�I ��A�'��A��5r}���#g?U����b"��}@k@y��T
פ�o5�q��lq��^؍���f�zB���yk����˽��}@ۅ�δ�γB9$m�jP>)W�d���[�fNd}ui�O}�Ӯ�w=?%�*�ސ���l�G��u�<���,D;ɲ�1�^�e�{{z^7��_�h�jH��S��:�w���y�b��X`\`�9$e�äQ���n=�:&�Aޚ��{��J���"���J:?d���	�f.�梪 �<F���������󢪍� &F����82��� b��f���j�˂�*�e�Ŋ�q��1�����R�c��/-���5��kb��9�x
[�|�&F%�|��O�Խ����	>��I�+���E^F
s��(~W�!�9s��U�<�Ua�lM�[�֮4��:�SΘm˖o�L���-Rޝ���ۆ���%T,��{�ֶC�ٿ�,��bL<�P�d���r�(F#�&>G��O�8�� j!;�9Nw��;==��}a�����q��G-�ݯ�h�l3a�S���	,��ކ��U��D�z{�[_�u��Xww��#��-��v/�ݢf.���cD��⎁����5۠�/���2���]��ϻ5�A�hJy���Ϙ�8.��sw^���<	�r\��0�j����� {�(�r-c[Mdؗ�p�x'�cK�/V=�\��U�f?ߑ�����:ߋ#�~� �[��o�?��:Q��|�]x�9v���Z����x����>c�M�6߲��4N�B������s*����v��_}�
Q������K�+�K�bj�=*3S/�74���TOp��_��� �#�8,	ύ��~�Gp�Qd�);W�
c�KcA�Ť�����H=�X�i���f/�L[8�QjU�L������9m���#�왡�`T�v����?a�_=�cq׃?�E@I!ۡ��~�; %�q�ō���
Ń��lT�)���u�b1��(v���B�*�5J^T/�"�����!�W�R�;*�W)��Iu�D ��y~G�I��\�ߓ���������S6��a�
۰�\�T,���Ӻ�h�����V�m�}��P%���뱱Z�z�����?�s/��s�e$*�������Y��Kp��8��:y[���~M<�8#��u��~�7��O�	����?/��	�	��9y��M�ădo��*����:�8dmx�#}be��4:�V+)��l2d����0�Z��]���W�VP��?�\/]�����ON]�z�5M=�C숚0d�:hᡂX�
�dT�w��'?�I��_UQ�i�"�KZJ-@��2b|J�L�d�q��|Ϣ��,>��1�@U�gScP��XD���Ăǵ��S�d��x�������[����U+��mݚ��s��a"Q��W�	/�R��m℩v�K^扑P?(�<W���Я�q���J*��� ����<s� )|FYw=#�-C���Q^G0>��"8�;n����Qi��_��
�ؓ���xl����Rɪ�U ��B�8��� `��j��J�L��R��j%�V󖌺a�g2m�f�����l�R1���^�(8c���	�����>�B��,jh�C��G=�g\�DH��Ģ3�yM�9s�G?��� ��t��\��e؇r�xxT�e�����g�{�g(���8 ���F�-�	E�ꇅd0�?$v�����im����4�q��\gϜ�
�� �TUO���&V��m͹Km��gӧ�ɚ�g0���\��,Y��ZjF 8����[���|�;߶� �er����Ӟ�v�~G�GGY'�.�8��<�>����0����N�~�wo���O�濽���|�K�Ї(�@������Z[�ڑ�W���;��L��R�y�ZD���D3Ed�{�1 ?g�֘IX�4�HH�'R���ޢ=��6�Xƕ�R�-Yl�����Β�����&�#g�� /T6/�.�'W.�A�( ��Ή:��/2QJ%3�<}j�6���>�5��h��泟�ĳ�	�B���'@�<�*����8@�)>`�J��liJ?s�|��͟��,Z�9ǎ���-Y��ҍ��:	�C� ��c�P�͚��s��k ��j�����p�;k��P�V��,�t.��۝v�����~D��'��'���=P���l��[-z��x��>�/��)��܋�BA�u��[&��� �L����+7o�VOo���|�V��54f,ח�j�&��uM'3�
��i��fuB�����ِXLLJE��sTkE��+�<U*T��x�6����'��9f���V)�)`Ԝ�,W�)�,NF �A-n�.��s�vq�S|���:$9Tp���r�)J�׬d�_Mh�տ* F�H� �s��l���7Nd)��T^	�C�|�!���`��}��c�(���7��M�|�9�dYTH.���Ch�hu�W��NU攬��J��C�������?�����"+�������k�xUO,�Pճ��[�f?@���V)3��r������M�5T��S�[n��ٌ?��ɤ�ko�굽h����\�/u��� ���}�S���� ��5G<_.xŀr��� �΢LǼ��;�rȪU����`(I�ChH3�紶�GO�%��j^��R �d<e�]�R�;g͚��D�]R���b����� <���pl���冻����RkA&�5���C=�t"�T��;����l�\o�%1KE�Y��L���~���4�f�'l޼C5R�����I^����=�3������>��Ɉ�x�_}��սB%�i��JU�D*�ႊ/Z�e��y�O<���a�w��.6 Q�3���M�8��А�_)�d�B}�������F�-�xy�{�;$��PB� ��Y.�Г�8�k�
�˸Vj�qȠ`,O�:���s��	���P#��ڄ	Y;c�xKF�J�B��b%���[`/{��f�z�X
��q&�F����t� ���T&��	�x0ڔנX�EmK�Y�P�!es�Rq�l;�앎3fd�!���7`;w����l6m�R��r}��~#Nk�r˖Q���p��usή����y����'O����ϼ�C�����(����i���z�������D��FI^���5�k$��'|�l{vo��{�ZB�M9����T�|f�>{��m��M㖬��;g�-Z�0���b$����M�uY�xp��p�yNyB��ū�>/�	8������s��P�����ࣨDIe���ܵ���n鲅������;�UvA9c�����[�h$,S�%X�x��G>2T �kW�k;�:�Cc�{Q�,�(��w��]�HhA#>k�[�p~���퓌�N^_Tm��œ%[y�"[�z�{�rɒ� �4aǘ�4i�m��+㖈g��o2jd�blE��찏�|�{|�����k��z1�H
ʜ��G4\}�r	.��R���mΜ�^��Z-{��kjj
yh>X`����8�U(���T9*�=� ;����ͷ�t��i$�-jw'�Y*�����W��[:2�r��^%�h�;����O%A�ep�t�'�����A4iy�������+eȜ�J�����^�:.���������'��6�f� )��2��Fk9p���!���[&KY�͝7�� �.X5�s����������n�C�!X��5�d��A^4��;�6���+�:E����=`-�d���J��������c���a�(XI�h��D�W�,U;�Ia�����իz?�C�� �9�K,W΁�c:�V�7d�3�Pq>-Ķ��\%OX�Tϟ�>sf���z��r��֯[i]�֬�w�'�(�X� 64N��7\��o��P�Y�3��vx��ԧl0?���^L���8�X�'`�G4�(-l��+^��v�K/�d�R,dq����~2�T��=r=�rr���1=��\!gY�Y��?�W]��+��=o1�KE��)o�r��+�寸�z��z��c�;���O?��4M���sV���o�q&{���R��LQ;��XT
�s�Ԁ?�1Oaokuݶt�X������;P��С�ֲ�U���(nc�ۻ�m��O*M ��<���#p	�U���e�SٝJ�g0�z+d�X$FRA��x�3�:�S@ �PGG��h�W�,��� ��w��k��G=�K��:(�DUZ�	�sϪxn��f� :�?��O|���:������+�Я���b�@f���y�{���.��8 j%Ā?qU�9�S���D'�@�b��X�{�!����q[��L۸q�����W=�Z�ĬTIZ���I����.�rm?}|�ޛt�-�,�RZ�����+(m����K/���Z���ډͰp1Wd$�w��K.��z�o���J���ჶ{�km=d{����x�2[�t�-X�ĦN�IPK�����py���S���:�����v$�'��I��5kV�u׾��zl\cʛ��w��F�L��'��JO�\�
%���앶x�
�\H�ԜEY�L`$Ȑ���CC�[n�ś8��-o�^��eM`�SO��H�hW��9ܺϊ�ǭ����./�J5���mv���Ya��/���m��%6�l�Jb	��4�*p�:!����� rq喳���LX���G������f<�A�99�+��h
�!��{��?�f{G�, 	��$� x�y��\�V����Զ'}�R���BQ3$�\=��0d��/@H	
��P�;�g[>�}�˸b�q}����%m6c���|O�H�J%)��kk׮���W�%9+�l�3�-�Lv��3M6c�\,Z�`p,�^�i� ?���t�v�H{�;���hx)\���h��s�])�':�wB<d��q��gv��n��ͪEK7d�!��\>����	S�׮x�M�1�E���Wo��:;)�w*˿Z�>u���e���-�����s�H�IC��7�卶t�|ˤ��Ҽ�J圵j���nO��S"��.Y��{,W0L�;���>�$�Pޕ�����?��ݪbB�!�]�U|��x�r&&ނ,�z����h\�l"c�Z�b�۳o�:�-I]F�������m0t�( �9�C��e���^|-
�LLx\]^
�62��    IDAT)�~>��[^��ƌ�� 2H=�(� {���3^X��,7�|�?T,�_� cE�)�鱦q���0��Sr�cqn�	 �o.�.�?��<lG2�T;�6~�lG�K�$rn	*�RK��@�cɰ��Nr��^�YI^!˶��$��D���3g�V-�������Oٔ)Sfۜ�l��Y�;��К��\�`�����B���s}��G}�p�Ϛ��$Ç8���L(�{���X�R��Zﳖ�v����k�X�\�*�:��*��3`�J�~�^ms��̦bw|�{���ĩ��-�jq��iם�U=7o�bOo����}�M�b���7ؔIM�L���߿��\��K&:�<�-&D���6�׬�Xɮ���p�&����ʇ����qH�-��ʾ��/����E�B&�it�gܬ�kZ��l�� ]@��a���Y�<��Fk����1���@��X"fK�-�ӧX�B�PO|4�_*�MLZx]�E�� �	��k��?@C*�1�O �!���W�@�<C!z������\<���, �&���/�=���|q(��3��L�c����;��qh
�V�����".�^J5z�b���s}�A�ߡ��XCn�)����e��"2v$�4�<�-�)���騼�WC�
���r�f�2���s�F"d<��Y��L���<��-_��E�]���"�z�s�>������&���?q�,��' ��w�.��?�q��p�)X���m{�^K���>|�r�3 ���í�֟+��`ͮ��7m�y-��؃?}�n���!I�H#,j�~����+����{ð�O8�lz�2{���n�b�Y�h�����K.���B�k��:�&����m�uX�����}�h�
w�x�j��B3��Q3������2���Y|�!��1X̸��h� ���Qy�ᥞqK[��ʃ�M��%����`��R�X��w�p-��%K��i��Z�I$#�?��kf�cyj1�u� �[Dfn��H��ol��'��d|1f	��H.[� ��6xdu��c�d�m��$��.ՖȌe���� �l��N W	d=�U`��9����A�qY8(E���������op�d�K3Ͻ{eT�_����F��T�_�تs�؅���E�Vڂ%묯��|��QD�0�jV3J��	ć�|������
���44��ʜ��	p�k,d�Y ����v���k������w�[�l���h�-���<{��W�kw���nhN�6׮�������<������7�w�g%*p�G�X-��,^do���J9gG:�O���]t�:ˤc�ܼϺ����N5Z{{��,�h{���k/p���!���Sn!/��c1`v����,g^��s	(U��p�O%_��q)�{l_�6;ұכ��h41n���y���	�Ƭ\�[�Ry��5�KU�$����j-�&$�- �1��/n�I���ǳTޅ��#�@��ի�k �xW�?���G��]%�i!����'�!�?5�1t�E�w�=�`_��j��,V|ǘ��e�3 #���^ƍ(%�˼`�S������v;��ɤV)����K��ɂ�x3h�E��;�S*�J�l�������
R�[�\�_�xc �Z������#�g��'/�6�������@E<)��]��kw���v��sl�����������;h;w�l�dk=|�*��}�C��K|�o>c{�����ؕ�Y��)U.����J�~;��a��/�`/\g�B�;��	L��%����n���m��|�*��UW�}�{ߐBCV>3�f�r�X8X>߾�;���HT�� ���p2��|�FI�����юfk��g��#8U.��4Xs�ѡ�/��ր�,/ i�W��(	�[t~BC�09�������H#�?������L� `�2� fx}������E���w˾�U�vޥ�����{}�R�����'s��{?��@/�P �ԩ��`,b�
�]�{M!�
Y4���!�,����ˁNT�<��Py�(���o"^�b��֭;�6]��9�|+����ON�e�W�5�ĳKZ*�`�\�
v�P���'>����V�<ө7����@"��C���K�Ƶ1���b�o�������s�^lS�N����T��d!_��{Z�\IX�^�TR�я��������ܼ�KL(��>��l�o'��e�L�2�>��?�Rq�R���v�7l��U�y��փ^���?�tο����Ÿ�i9f�6]����kM@V�5�U7���7�n��@D�`yPPj��[Ա�57?cm���ԓ�.�(Y�"�Z$i;p��ԓ ����A�|*�'�%Ǌ��U@˟=E#���(����� �����qw>���ƫ�3�/e��r�ԱFh@���>���fl�p�, +`��z����?� �j�����[�@
G��)����˳y��}�f�6@kB�
�#��sqN5p�����4~J�gSc�����V�E�y�ԓ��J-m�M��i�d;���V(�,fiK$�<���ϸR�8������7W������%�Ur��ϝE<�tv���?�|�\k�fl���n8�����\�v��o�x֎w،Y���kǛ���:p��-��8O�����n��m�}���߾�ە�7���皑�>h�����h�_�-�?�j��=��}6�����`_xў�D���l9h�����]w]�����C�#���G��d��gR�s&�{��׹��-�?,(	8�H%���쩧���foW�M'���Ja��	z�v���<hǻ����=���z��8��8QG��:	�"Їw*�s#�`� :�Dy��~���=	EX�H/���*�ޱ�6�S d��R��&���]���O�'�:��O7.���E��wj5�1X$X��s P�]��(s���i�GM�J%cV��_{�'yŬ`U�7$wR�N��K_a�Z��unt�X��ڇ�\�Go��3qy.h x��_�5b)�7�����~N��G�w�0�bǺ�Q[T`qj=�i�]��~���k�`�7\�E�ܺ;��o<'�o�A�?}��n���[N?��r������e$��lX���]�Mv�k_k}�]� h�mmV*Z&s�����~/�0q����W�����V(E���o�;n6�~Ǫ�A�U�� �.#:a���z���E��re����b��sO!1e����b�<��-*b&̛� ��%�p�r�#���)��U����*E��$Y�����g�i8�
t�/�MI� �(�>@�"�o��+I^�Y$��*����0N����2FQ��v�w��E���)�E����N�`'�㆘eh<�c>@��!p^<%��1^��s�Z�	w,Q���Zb�֞c�t�*ł%��n��9e�6s�W�T+�ư�Qǅ�8���˾���9�so�L�ʰ�s�����S�#۰�bPʥ�#v��>��hsj���R%����H5X�T�;�Y2�`�����S�{ىo~�[�ӟ>4��)�v�������t�y$�@�/�\qk捿�z�3w�M�`--{m�Χ�ۭ��{(U�K�Y�m�s-�j�����N��Kd3 x�b�o�8��������@F�dU+<�QGh�^v�*�56em|R��%"���$���Y�N��Q�ki�|2|�zEQ�ꑤ��3��=�p����τ�?��Á?�*�1h��-����1E���0��'��z�� ٗE�W�I��%����3�n���߹�[N�`�(X,%��������@[��)��?�#��8��L���;�4*�2�K
�z;�9�ς���ȅ�&Mj��&{UO/�Xt*��05����T&�4Y���c�]In0���Ɛ����3���:���-���	�f���Rgh\6iG:Z�8���;�����^8C=�����%�^fM�B������/���	���- ���mw�z�WO?���>^ځ�?��^�y筱�_�?��?���zmǎ�]�s��O��d�̚� �R̃��H��%��ÝE����o}k��?�4z����?��?��L&ܠ�����?\�77�k��X�T�$��(Z��)�ʖ�d�>�%�F�^������j�Q����_��M�ZU%�>
62�Ƥ�?������v�n�±������^x?P����{
��E� +@�g�ƍC�d��J`c1�P�*���n���;h#�9 �𦼁<Z����������Ϙq��ba9C�2W 9�sB�: |����I%�CU�t*���>������:}W�%~=.�%K�yrd� �<�RԎ�gt��a��_�eμپ�>��%ܻ!��c�!ཽ���y�HZD=zĽ�'�|��Cpl�˯Y���=w�M�8œL)�����ǝ���t=aQ�$�1�$M
�8���T�/�d��f�&M�	��Z|����n��
�H�����>ॺ8r��ċb03�xXE�_�YX�d��
ϯ���`��m�3��b��~�R����
�Wl�S;�)�b��*D�����$��(�� I�	񏴃�B��`5�� {��6��O@�Z@Ř�l����h�js9o�5�v�\�9- �D�
�R��*�'ޞ�]��Ї>�/Zs>��Cm�c<��p�,
@ �x��P�?�$I�i�H�/c
��j$�
�k�܇J���Ϟ17�}�'qkkk?��1i��?g�$[�p�UJ�fR�P�͛�{����W���L�T�L���.X�Qt-�W�5&Bc�8��x2�B���/�`	�=�1O$��MQ���\�%j<�����$�
100�`WO�3�|X�K���7�s������-�e3Pqu	� {�ej��w:�,2q,fl+��Fݐ��=�)4�*U���X;z&��%����ޡV�];�c��<�Db
@R�/�g�a{��^���>��͎���9O����
p���ͽ��[�'���;T5��0��?���ͻ'Y D��0�G<3���w��|�� 8�� ˛y�1�'��Up�xrP�Gq<��}�W��@P���W�wE�n��ÜQ�"2��:��Mg@s�>G�mBL�RW�y8��k|�6h�Zf�_mF�R�X"��$ǁ���k�lm�Ԭ��B	�Z��嚢��2��_�����Qo�y}��/�o�>扏0���
/H
 ����3\��c`NJA�*�2Hهg�������JMwZ���-������Ƒ�J<�1Ȕ.���dnP&/������->�^kؓ��2�M�'��ŢW�� �%�TUO��F����3+ێg���P*��Y&��~�P���Q/�Lc5���._�$<Y��OF���k��^|X���\7�/W&E�d���y��7������ċ�nx��HOJ�y���&y%t%�_�+�|��R���U�Y'=� 0���1��X�(�THF��J�
Us�1$�Bu�6� |�L�W*��E�%�W}!�����چ,�����β��g�b>��wN���Ujq7�[{�7�
�@������y<^�Q,:<G����s���<&�8���Y��>�яz��W�A�<+B<8�����3��𼠿XP�����d�c�?
F�
�UISJ)%���jG��s*���ZH���AY�|��h�نA�W@�Z�u�	��*�'��Xaox���4�8ٵ;ةZWW���{z:��U:��������w�O�y��b��-^��fϙZ�UF���LV=i�%'T"�\�z�y��' �V�, ȭϺ�������"eч��pT�$8q (G@� c%�L>�ˈ#0�⃪�0��4�G���ƈ
�i�H&�W�.�"���o|�ϋ�EP`9]ŠU��/�|^�W�7��%�CUφlҊyJ�������Z]�>V1yz�O�4�Θ:�/^:y�)�q��>$-66f=��2����н��w�*j')9��j� �澸O����IU�ERυg� .�=F�:��^��H
���P��JӧN��4�z���K@%i#��˲R�h���|��>�C��,��n��i!�K�Ë��L�b�xSVw4�cB�`�H�y���\*�-V+Z__�<�ú�[-�E�@�Ѥ:�e?��a��H����-�g�fOwz(^K�j�s��X5xUp��&`�*�� դ?�e��A����eA,�n�
���$�D�;�� ���Bg����{�2/�`̊Ҕg��\΍�1������,M
����;D���3��x%|8��Ca�V�N^�U=U�٬X����t�rܪ��%bY�5�L�4y�54��L��
%4��~PBC�[Ro<ݛo�Kf�ӷ��Z�0i�'�a���H���ûG����_�Ǭ���L���^f��,m%~1�����j����������#�<|�i�Ղ ��� �@�`��~y���$��!@�Ń�G�n3����眀?n#�q��[�qo�ސa ����Xs�6��h������;CU�\�b� ��ϵ9s�[ie���*�~Z�4�����;��k��P>����C�/�%�幊g,�D����AF��V�!N����ƽ��Z�%ٔU�1D����ǖ�,�EsPF�"���b�x6m�<T�M�ζ
rj���=Q��,OEU=CI��4%ɻ��ϱ��?Ǫ����9�;g�^`����Tz�W�-�V$^���{�*������O9��
������|�	�X�h�U�n�h;C�.�AϙsS�D���/�N����2�O��W���)e��B�W�/\�.^�"��Lhd�������Y˒���-�4�xMx=h�D��;����IKO�[oO������>�S��w����'��b�x谵t�"�3w�U������g�
xVr�5����+��|�O�J>�
���>��{��� HW?��g��ƶ ���q���b�y����U�K��~
��#/�G�D�Z�W�2�D%�k�˜k����Hj29�P=�J)�}NJ:��a���a�ٖL�Ӄ�l�|�*�:s���d�s����H� ��<����3_[�a���}th�s}����
��QZ�1�Ƚ@�To�K�g�g�©F:||���UKގ�������M�z���?EwM���������{��]������ٚm)�R�Bh�iIDEE@D=��S�v��;˝�������"-	M@J	%=�������g~����g��eg7!	p�/^����Oy��y+
/?��4[nHic�nt]j'��Uf5��aM�N9�\@�� w:@l:!k������+�d ��;�c��L˺\�@��ƣ�-EG�Yˮ���?bd�U��D��W�o_��&��q�1P���������\9�����K��AZ�\RH��z�=�G�,;eq�:��\~<֛�#���La�tMi�^���w5�rƿ�y��|7��9�����!˘�ƌ0m�1���H��4Ǝ��c&��D7�`"���L���η.>�hU��c���+ĭ@�����r�����%4�����+��!���z�o�Ĺ���_�O�s���b��kim�����g��_B����
�� �ߵ�\ʙ�d�b^K�T�F͞��c0}���$0��Lw�:y�N��G � `qa�{'�/�+��ͨ�9�#�X�~��e�ǳV"�g=��7n����n��O�lZ/|~�����C7�+��G?F�<�2�Hu�J�R��7o�|��	�.��8q���-��;����m�ē��r���g2�T�Z:t��7�+�c왑6b7�Dp��(�,����� �����u�x���0�F` ��4-2���T�沎���5��w�)�OO���D���`�UW]�g��>����زy�ݻ�ݽ����Ne՘�葿Z'�@0
zy�Aq�V�Z�Jf,��9��Q8ɿ*��/�3�F�Ў����-��M�g�-r�PUgvЏ�3��S1�e:1c���1�D!��.�E�4"V݈��&6�    IDAT1�(+���l�p<��+s�y��i޹RKU����,k��x����R.������P�/5p|�n�zj����+-_�kZ���埓�HDҚ��f��ڠ�!��Kn�~�ݐÆ���m�J�}�D
ȧ�uTU7`��Mx��g���ΰ-]�ʍ�EC)9����R|>��[�v�]mh^��څ�
_��&Rq�T'`nݺ�������E6݁3'�S���O��"/�;}A�
Q�3E44�⤙���u�+M)�ƸX���mZ&�=͖^�[ɋ  *|����O�'�F�P<D��4�!�/�2�����|�L�S����ez	��wU�������_T�qoLA�C��XA��Cy�K�����|%kS�2	���g�ƭV�L��9�I�X�v�Pd�����ӳ�z����,�s�F�P�@߱#?�k�a��V����g��������i��=���'��O�fl�(0��3��"��aX�p+�"
�(3�`+��n$q1K��\�$�:ȏ�y�6V��4o5�SXB` �oni�~p��/���3jk-2oZ�I�B���r��l�
�޹�<_ח�Gn%	 Å�@/K�)������?�ً�h !���2�Y�C����6nي'�z��$Ba���p���1f�XdҎ(�ii,ء�G�
��:}h��v�Џi15*�����ػ7n�?ӧ��I��ǍǉӧXrD8��c*r��,�ٜz��5��+����c�f(ȇ�A��`v����H�6��x ^/^�{����'YR:KTV�>PПn�A����+e�w�V~6.,C�)3%�W1
�L4��*�#)�;p,3RE;��s"{��2�'p�e�_�p�u1�U��#�w��|���j$��رk7�T�Y�R`�Xv�:
�T�hXiL9��<��޹ۇt]lh�c�W?"!Ge�HvPkl���k�oτ@����$��#hjn@.������ѳ�s驝�Rɜ�|(���'];Ѩ#g����`��b?^��!JQ���tv5D�Λ�"W���4�
#p�e����"/i�^
N��i���J[J`e��xj�fJ��o���6y�
�tM�k�tHiJ�R���S)~��?)����N&��N�F�
WYos[�� �H!V"���#hjj���G�豣1��s0bD�-b�&�@G�������7~S`�����%1O�����r�e�oP>eA^��ٜ�1�Ҏn�����|��cu�ً�Q�8sYa[�q�- ���:
� � >�w�gT����}O�K�\b	�D��*{/�����`���x�����N��[
W&�᭭8��3��:�t��+-�i`X6L��u$n�D�P��ތ!	����{L�����a@�]]��gFO�˸ TU$�t�?\L)�"4o�SE:����k�{fΘn)r
R�`��,Z���v�!��"+��O��%�,K�x�����%ȿX阞�;R;��[�>�j��x�K�;�t�"38x��딿�wޏ�+��5��3��Vz�W_w��������RN��}l��4����Ǿ�ml�Ej�|�|i*Ϣާ�x�/���ۘ��|�����t��c<s{�g]�[��7��,�h�z�����wߋb!`����(��DCat'2�j����t�"�[�]��j�c����k��I�����5�� 8��;X<��q���G	���~N����>��!�����b�ݟE^�-�7J��܋L�t�����(䄾�k0m�q�1P�3��}o�ހM^���b-�T������|ģ��r�x}��e�9���(��ln���<�1�&q%���D����5�*�����{����ꫯ�s�������h-��4���f@2�s�������o,J>�6��������]>�t��b3�ѕ��3N�[=�'uD >��7(��u1h�̸#D�~��]3o~`�!��?l�� P(&m3�Ǎ&R1����#9ʡ�;��H#�A��n���Q�,��:�*<O�ŏb!_ dϗ�q���E����X�
pj����ek��Ϗ"��C�_4�y�	���2W�sW���S���Q��A�g��@��5*�2�.�r��vr�}�qN�
�f��h7?n�
șu����}d��d���B
���(�Jb�I
�5k��?]��_˥oz��t_ݟ�{��ʲeϛO���G��$`�u���<�����������u�7p�N�gL���^ U��woL�g��{Nq���8��_@??c�n��P���TWע;���K�3�i�%@K��>AG���5҃��?��������\����p���"��D0����²�F�le�y���	3����)S1|�([l�,�]�|�M
?�{��Pr����j��U%�O~�S��\ ��4P���'ٙ
*�i[���Ի`D~CUHrQ�r���]XR��~_+�+R+�
sA�cˋ�H&�6�Q�E�y f.8���,V/P0.j�N���Q��[��aaN��l��,'��;>��ʆ7��;>�}j����̆�.Y�
l6��X�h�)�%���6z(2�iS�dQ���&P��p�B��}���s��2�>���RiLl1�$`��������i��tPd!R>ւ�|V��/WcB���B1�N�0���=8ͱ�w���~nŜ�)�.�bP���kɕ�ci�X<���_����w�{�:��c	jn�l�*d�7��dZ5}Y�
���W�p̵_��A�We�]����u�x`*~׻�X���	��.{o(&�z ��^���fR���O௩�K9���w���a��عk��SScƏ���3N�~�������sK���O������:�ނy?��;n���,���8G�>��C���LC۲e�|�Q�;���0�����ο�ǉ3Nø�l�R@��G?*7s (35졇�x��i_�U>w�\9�L�,�O�� %�kA{ϯ�a5�8��6H�Ks����ٳվ��B*܆�a����5��!g-n �Ԇ��#	
�S{$�dm�>ט��:�l|SH r��M;��A;߹-r(�]@�.��.�Ի��&
�a�%����	rL�%�����/?r)���!�r-q|d�p,,�C?p0�xe
E
K�E�\|��ˢ�,�Hԏ|��K�_��~��s`��Y9� >Q�	U~���06W�sI:�Ɓ�E&�:�����
~�r�oB�ד
�s~ow������(���|�w�C�	�r-վ�/A!�GkQ�@�W�C��*��Ԟ�P9u�)Fa�����Q�����2�g�����g���n��I�Mwa붍xq�2�]�Y�c-��s�4kƑG���M�X]$���7��'�3}5��_0�����gZ��ITǪp���ٳ�J'��Վ�;6a�ڕ�XҜ%v����ޑDC����ך�g����g�d�YH3�.!���z �+'����ȇ��\���'��``��kj�Vֿ�x���M��9��,�ȣ������hf&����ȕ���g�,ɥ$�1A��1wF �l΁-�P0Rr�el3�	v��c	�sHf҈	�A��	������cڤ ��|�H0T�hx�Q d�����~ݿ$t|�����YՏ*ӈ�'��I�܉hU�	��6|���m�Fb�:��Y��C�e`�-����y}Z]�R�!��v���>��6�����|_�o�~:>G՜-�.����.}���o�G�����/o~(ʆ�xȚ���ۓ��������X�E�l
��*g�����4˂+Q�H����)�bj-���B��/�Ӂ��ͣ���ǐ�¢���g>��F�F��R5Y)Oz�����>S>?���5e>�B.G���ذn��چ*r�\&�5��b���v�L�s�F�Θ�/�+��)=Ͼ���1�����ߏw�o���S�rݼj����$��a4�U�ww�S��d"���6��&����۶�D2�Î])\r�[q�Ygوs�٨�����G$p���[���Z;"�Y ��w���hCie�@�/ ��UN����t����H�ՍƦZD��X~n�u����[�)u�+~�3��O],�@Е�s��s�s��;���Q����(Z��I'�� �pO�����\�֚�F��Ӊd"��a���]�W@�#Lh�K&��8] 4�0���sYz�z���6�;�C�lٺ�R[Z�͔D?���_&ldb<���	�g*�A$\���v�wU�0������%�3�``n!]
9���v���)�ڣ��khmѰ�P������u���;�mn5���F��b$�j�N���o��xI(Ïp��d�w�Ecc���e�0Ǎ�fKZ?���\�,�0v��_ l���xD�Ae%E)�Rp�n�Z?X�_�Ϸ��(��8��5Z4	>7��I'��/����g?kV�R��\<��<r�n��ғ�2��y�F��1���-�͛v"ѝFWg�]~f�<�((�)��寑+d�)B�m�q�n�_�����U_!h��Q�F�s�������v�0��S���ֶ��7�`��lټ�`5V�ۍ�Ǟ��~��f����]�(���G>�[lq�zR(�˿��� >����~��D*gn\o��P�}�9�����|s�<'�e�П�!�u>��[�@�B۷�㩿����{pͻ�j�'���R�r�_je��H����K�੿>�a��8��3Q[C��TbOp)�-L�n����~[6n�I�gb��1�{b_�B���{�X��R˪�d�YhF��T9�aAD����]���>�V��g�Css#�:�4C�
`�8�A:�3Mه4�LWdp�
�x��'�Pi⤣q���/cq(���A��OR� �q[ :;�x�'�Λ;��KY#ΏO!@߹��KMxؐ���������SO��L���5wV�*��P���}x~�Kv��SN��)cM ��a�@�IQ�_)S.��aǮ��랽����X<����8��	���o���;z?,����5F�C���s}�k_���>����Y�ϦM<�^����FMT��ɿ�c�D;���?b��ᨭ�F�Ƶ���0���JᕗW!k@[�5v>�w��^�;v첖�[�mvsPR�z5��_0�{������E��TL8f<>����V�Z�g��N<a��v�؆T�u��ՙD[�&���qL�|<>������I���B!S&ӹ����'�P0����C�Z���Be���J�/]��WҾ��M�.-���@��-"�9�~��Im�\6��/��IG �ڃb.m�j_>l�`A�b�B�y�`;vv��G�!���/��p��@�im�&�F�`�|h2S���kVo�#�=�au�p�[/E>w�}�8�R>f�d���?��#X���q��:�(�3=�{�=��.��L*��}��q\�΋P]4�`UU�4g��JUz�e_۷����?��#G��K�"_ �e-�)�r�&�g9dr��b@�����59n��v�t$��P`��#닙h08ZL�62�B��r���9gOGsK����Dssn�S*��*I>G�y�V�}ϟp�)'cƌL1��ǥ�z}�.5�M!�!��%�-�O<�3�:S���v H� A?_�b*�|ϴ��c��v,Z�8�	��yfS#�Z\����^% � �� +����-1� �����d	�%��#F��v�l��n^��L����-Ƨ����OE��?kּ�'�N�6MMðr�ˮ��AgWk�lB&�N|�����_Cu���.������+ʬ�ڻ�̟!���>Ǖ}��q���o4M�ޭ��Ow��9�M�ݲ��DW��#�Ύ֭k3�߰1�	��7-^��� ��M�� ����ċ;� � ��A�3!�23�߁}��\���Ո�ʄ���_�/�8��Y�8�� ��c<D���M�C0�3�~[�ua�%Ȥ�����Q��ȹwf:�e��4Sr�(׬m�c�=���:̟w1�$KrJ�����ӓF��j<��X�b5��9�?�l�U{�h�tG������,��YtttᲷ���z�I�O*�	�ְ���lX�>�c��/:��=�D�˅�D2�@$
�$�r�0��V<��X�v=��0	g�5��N��R�9b��~?��\���6�����~�aÚpڜ��:�� �RK��y�Ɲ��_1>�c6mڂ����8�sp��Lw�Ͼ/��K��{'��!�z,_�
�?��<�TL;a<ry���A��qə��4��wo
-z��.k=
��rZA�V��>�����Q�>�W�J%�����X)ۇ��~T�W�5�D��/Z[M�a;����wYV��X/�y�[�����N�3@W��5+���s��!d3�\��l ]�Y��E|埾�`�ʺ����?�굫LY�{�/�������@d���#F��|��e\��n��4�8 ����TPƢ����[�+D�qs��x
n��F����n/�2������6,\��x����9g��{�5��m�L+@���[�l���c�+8?�@)n�]���Z�3�8�=g6��X,�7��#�4ͬ�1�7RÆ�Y�ޓ£���T2��_~b�r�����ϥ�Q2߶T+^Y���|��:\�ˬ�]u. O͛�T
�]J��F��ú�m�5�$?}�{}�s'���'�s�JK>C|o����i\z�h���=�����/C6�|�e�h۰�-�*��r��"�NWe�u�.����g�o7���X��q�_�f.�c��|�k�1�KQ�b1��N��f:+5�?���w���0�1�r�-K�.'
�_v�"	 �>֮Y�|��~�N�Z��;����Rx�o�G�2�=�|�
K��h�������cǘ_��DP�G�>�y�|��?Sx���ٓ��E�ބ�e0��;�̨W����װ�����J�+�{*��
��J�KqM�'�?�f�2w�ҥK�eFk��t٩����i����	ذa�~�^�7�����/ K~.�zC�wc��G�c[5����'>���aX�n#~{�-�M���R��b�����A��e �`J�>������z��]x���8rT���]�{M������љ�捛�i��j/����5r�Pkb^��f�?>^y�#l���W��c�a��ٸ��������M �8L�
�-i�}��p���bx��U��3�.�ɓ�@0�u�UV.����o �?ņ�x�ѥ�z�;.B4l��������X�ڳӹ(~0E�P����.A(\�K.��/�p���L��.64<�ebVK��۫�x�_�~�F��'Ok���"M"/�P[_�\&��D���5�"�L��������s�%� VC-�Yg�nT�� ��a�0RE��*{��X���3;����ٵ˄K0A6�<�����ۑ�&QS]o.��x�<�֬^�Y��a��V���teutbյ��l7������*��;���=6�����OPW?��2�v�4����~��]���?`ƌ�s�$:��]�1���z�5$)+��T�a�O��4������ǌBw��(��6!���+�D��h�hG
�0v�N��+���E.�L(�]q_��G�sޥ��@�k�B��ʖ7[HnQ���������R;ŧ�=̿�׮]kץ��Һ�3�O}]�~�>�.��`ێ-�%M7�ջ�CX��{�ص���}�1���Z�v�e����^�=o��/5J3�|>\r�[p�y� �����e�b������2��>�5u���@ۖ����_�N���~��X掸��կb���fR�8����$��1����shp�H�e��.�/ҫ����`��-XH��gҤ1Ȧ]Jlk��6����G�Y��w�!W̠:V��;�X��Id3�u�y�U�H�hEZ��Z1z�K�?�^�;�	�PUU��k���Ï���W]�6�	�|Y�=b�}�Q�ݳq�F�m���mZT8T���[�5k�aΙ�b��#-x�L ��Mhmn�豣-��qs6nX_���~�b��O��@����CJ8A���    IDAT�������l��=;�m�f�X��b�Mx��'��P�K.���_,�b�w��13z��֯{�V�������I�m؄�'LŌ����k���c�����Ƙb�q����B(�@���������a�Y3��\gV�)�5c��񨮪Ǯ]۱e�Z���.�T�~�I1k��Y�`ֵ�y�9��˦����-��=Q��]V���Ą�c�򣻫Ú��6��@g�[�m�Ν��L'	נ=��,B<�,k�ƛS*D�AyU�W���ڂ��H����}����?|_i��!�s�e���[�j�^V��|��!�
N?�t�T�g:�n�Kصs��@���Hg3�ҫ�fV�K/�6���W����܉��.,\�PO�Y���P�oni��������1�A��uj����x�ϓ���ш�n� ���ȫ=��>�4^X��Ip"���>� N�}:&N>U�l����I+A�L�d03D���>6u��0b�H�[�� h@����ޟ\DFJ��~>ܜX�:m�����X��l���w�-s���I��M��L<u�����8ַ����]����)�w�"��_�֋�P��a��5b�䩨�kp�7�70f�<�ϊWV�i�}�jq��������Ǝ3�j��Tr�Y�ʺ��I�i�},��U�0��,;)[�"�ǔ��[u'��\N�֬Ya��-�:;�x聧lc�����\�8��駝�|�o�[ca�%��3O����m�_�����!�O�=Z�����Fw"oEl�\�����+m�؋a��Eذn=fΚ��'M7৛�����8�����b):�v#��Buu=~��[��쬳g�e�0d30�9u��o��@8��ӆ�<i�Z���W�5n���'L7Z�L>�qG���e�3Q�*ڸa-6o]i� �b/,{�=�8�;�\L�t����Ģ�8y*��u.���GWW�7;:��ol.|�l����c�1ۗ�1�_�ֳ��c�o��,)b^k��\KS�Y����T\��ϸ�<�v*�&����F��شq=�a	6mjC!�A�u�˙�Hkw���8��3�٦r�=��w��]�v�ǧ��?����"���l�5uHuw�8���p�EZ��ݝX��9�̙����S�Zpgډ3�3���n�����ؼys��YY���������"�b�Y��O�w���\D��SS؟�}��I*Me����ތ �s�������QG�1�3���N9���
w�옝ǚ�+L㣏���E�6��[�z	jc�( �#F�ńc�������*dy�]���=F����ex������dc˴A�-��`�6ړD%ScGb/���æI�U7�~���u�}�Id#�5���N2_��9f�6+W���V��Dx���gA̿�\��ģ"N:�TD���,hcЕDy��6�>��ۆ����g�Gĳi��@um���#�M�,_�ľ�Фe�K/c�ɳp�qS-B��ة���[���֬{ъ�BA����n�bU8�hh"wL#F�������+���M'���{v�et�btIΜ9�O8��+hI� qԨ#��A�H8�]�����9 ��^Y�Gys,�j2��4Z��q��i���?B.��/����L(�^��>�{v�j���z�`���_��_���Z�5n��3���֯ ��?�9ۧ�����I�?+������bP����n�E*k֬r�D��{��ZP��9s�c���1�-��H$q��oǣ�>�)�Km��A��@�@>��?v�����;�\ǟR*n!�15 ��ј-�Ԁ;w�4ʆ�^z��wS..��'L�����7e���5�QV
NБ/Q!�����ӹZ��)!3��4o��g��|s瞅Y3N,q��L�oji��ˏ��V%�k�V�?����Y�=�l=�HG��Bc�(TU�ώ���S(����c1m7�{���G�Ōf��u����BC�00W���8R(sh߻�,��K^�Ë�9���̓���n��I4Է���,1��Mw�5�hߍ��^k�I@۾5�+��#��3�c?u���kh1����WU��u[����2�}̽�|�9�]{m\he�@2�t�w�EZ��oCw�?��ο�0a�DTW� ��Y�OK�&�
E�2L�d�;en#V���;�c[.�w	F��6�U8X���ᨎ58�K��H,׍ή=�h��K/��SO=m�o޼y���2¶P���Z˰���u�T�,���N��)�w�h۸��c�%f�dShj�Z�2;���YDcUH&��s��3	�}���a�fd�yK�e�?W����wߌ#������Be�y}��3%RhP�E�u��FL�"�Db��(����V�y睇�有h�4�R�o7� �G���R>I���Ltw㩿>a�E,2WR�׸�J������7���OM"��t�3�	J�?�S�֙��,���0�E��1N	ݨ��}��f�o,�Rր5����rQ0����9MEf�9��/e��g���(��L�C�|&n
ˮ�pՕW����@w�����K>Q�.�?�����"���M��M7b��H���e�����;j�Q�2�̾����sK�����_8��0�����d-��M3E.gi�N�8Ͷ�{���m�މ�-Ɨ��O�h�oFu55_f� ��U�1��&�Gx��'��_�����U��,!�\��L��0��-%0_�r���
��w?��O8��Ӎ��2_��1�ч`�u�rM;�&���g?�)V�Y���w-&M9�h�K�D��'��j*(X��	��꘽c&�ړ#F� �l�s�C,,еBM<C-�� 
�<>���z�U��{fO�n�,��9��S���4r��ձ�(���o`��Mx���c��wOյ5�˰��DB��,��*�4���;��o�4Z#�DM(H�z��yy����ތ�5��M��%���ܫ���-���ζ�<���x.����*c��!Z�sΞ��g�RBp�%����?T���1�F��G{�^hB��6���"��ń[r�z�5���T�~��@.�\�}�J��Hu'��@��#�iy��H�B]��n�fA�%K��ɕo^t�ܨ��\X��9������^z)���
�F�lق���[#��G���V�'`k�_����T�.����@�wް����ry\~����>�qJ��aʣ�8�'�p���6[�KKK�}�{1bdS)>�F����N�s��r���x啗��}����y�7o�c�$�u5+����L�|2���p����w[�ͧ?��3
���8��
8*
Z�Jv�>�X˖?�[n��=i|�_G��<�d(�ppEZ�7[�TM����p�w��{�ԩ���>`<F2jst�T�/�\�b������ ���obÆux���o-6	�|_'����	���eEV�`���}�߬0�C� �Zb�V��#���F,G�P$%C�����L%3֓��ʀ廮yg	 E]"��3��T�Θ�
�mNw�܍y�.��g�m��9����UE1˭�.|�_0��B|?Ο���[kwO/�����@� �G�2)OR����`���c	�7\w=�=�XK���c���5��Y�O���B���U[[o�>y�dL�t&M�d������L�,e���|�)l޲�h������
sO��7���6s鳙��L�&��<S�"�*�U'�{���䗮.�<�6,w��=V���=��w��]��f�� �3������q�@�[�8�>��{�\^��3��mWX���9�b�JI�GkJ��|7f8�}p�u�YIw�l��Vk�n�Oƍ�ϲ����o��/�%��s�W}�@��>��������+�.�m��vwZ��EpV���Kˍ�+�̚�B���j�g̜%��	aG����\�Ɍ�p��Ԟ%�պ��b�����������1���q��e���]�������|�Q�Z]���C�z(�'Y���*3o�k��S�rt����OBC6N��Hi�^0�k�87]ݝ��׿n�T�gS�S��"�ý��<^~ �oޗA]���7�lV(Ӻ�}*��r�������q�l>}.�G����ɬu� ��i.g�K�?:W�cj���|�u�p����-U�
�mQ�g��"���MWcN�?��?`Ŋ��;0q�D|�S��2m�iS�I��r�G=L�mj.Ϋ�~��x���ֳ�y�6І��o|Ê\�r:z���p��ӜB�*�a��͂\��R߄J������c�Y����3�\ݻ�F��X����.!��\Ι�Ȕ�}�=����fw��ח����	Ǣ���^承���5�	��ZR%�/p�W��SL���8{�7���\s>yi��p��'�ۇ
�2U*���;�k��`3�>[~WIx����S���]��z���>��h^��Ũ�A��aP�B���O��O��3œn^
5�mR0+�G�}�kMy�0SkC�$כ�޵��$ �����n�����������p�X������<����޻��x9�,��O�Q:���X��O~?��O��SO�F�R���9ܸ�ٕ������fk���ݍ�����J�����GW"� �]�����C�5�����0p!�s�y��>�7�s��Z��2��k�E���6��s��eQ�gq75�)U��[g��q����,S榛n*[w^��2}J\�|>+7�O�Ss��M�Vp���y���l�|^*�&�k��XI��k��(tLP��Ҝ�7�T|f��_ti��#KV��+i��%�3��?�߁������@��>��WZ��?Z����g̭C�g̎���ts�QY���s��ˊ�Kq�
Y�"y�>�?�'&X��N�﷍�~�Cop�?4��c5��4�}ьg�We�X�/�R�����4N��J��1�!^��z\�W_��JD�'�A�K.
�?�;Ǉ���$p]{��S`���ečB<���E4�p"ë4 �ݧ)N���}�ƍ+��qC����H��y�	��ɭ�}n�� �����bޗ�?��,i���:+Ҳ��$���
��j�^W�B�"AR)�J๪ %�����r���T��S�j���eM�	{^�;��	׃,!��[�x��i��)P�Q��?;����˕ƹR�W
��k����ה�s|��x�	k�Ƚa�%>�]�F���ԓf�U~dux��!���h�aY =-��&m�m����F$['9��`�� B��w�X�e!�}��ɟo��?�ϟ`Lp��T�s��I2���N���DN�����G���l�C!z��� ;P7[������U_U�����X�?�~��_ۦ%��%����njC͟�d�,�� .2�ļ����PY�CAI��c���3��4Tj�^�qf��`�K�}��Oa���,��֟���1.fi=��~��aM�XZ���������{���l�e��ɱ&s's�Y��:��)��b�.!�w~�N�JH��Y��_�u�[��������i��X�g8���?�b�0��H>����%U/�MB��� �<=���^ӫ����ͮ�+�Y�\���,t��(��뀚i���$�q�8�Y%*��1��]�a,���{��/~Ѵ4�T��Wr2�-G��[���	qik�*cD�A�=5�z�i�H
��n.��el��.����O�����e9h2t7�閠��?��Σ�e@� F0�Ї>�Oo�Jc��p'��y�FL%Gn����z!�݀�g�u�i<^�Z=�i�󹔦���5ſq�8�|g�>�@�8	2�Ko7��u貚z ^kDs�U<��z���޷T�{��������������$ؗ�X���:�O_2����4.
Uj�	�<N��?hr�?�k�߻�}B��]���]�8��N	�D�f�]�L��ޚ?��c�l+1��tKP�_J�/95p�ɾ�8���ÏW���ڠ��㩽3�[�L#R����I��k��V��S�3�ր����o��4L��ILŀ<0������7O<����]և��g���g�	c+�w�
����TO�+��FA�Ɨ�Qh0���)Gj�{��eE����_��=��y����j�e���d�p�6�;� �  -J�,еT]O���'MS8#�����/,p-y*���#����;��������.kS��ڽ7��w��˔���X  AN��Û�9�f��	��
�)�h��)��{z�!����� <� ����W�}�9�=�I�A	������[np
 �'��&�O�;��;��\��'�+��c$���}	� ��Z��b�6Xa�M���!��@�^�KS�'S>ǅk�V����/�嫴Β�q �+~�ؐ��v����x+��9�Z���)�%O�'!�w�6�h�Z���s ����pK�'ô!�D���+�Sօ6�ib%��-��e�-�|���8-N<���� @@��`/^ %ׁ�&z�M8������;�_�`����C'�D��Sȹ�G����0G�����	D�M
�@�a�����5���xǍ�4i�;�8N�|x�� �%Ùw����j��O�^vdJ�q������'��&L���H�Ф�4���Y�}h�|@#0�4\�+�b�=M|P:�,EU��v�.���T��J�r���6��L-���W�Cg�qo�NU�e�Τ'P3pK�?�2Y��L��1����5}Q�������a�)x�
�x�J��\�C=4C#``�(�}/�v� ���<NBA^�O��z]���zPk��R:����'Y�7ρ�Ţ8�9V� �	�B�-غu;�[�Ě�����M�''�Z�R�zg�ȊP�N�ƿs�9���|��ch��#P)���׊�oJɕ�/OS��3L`�8@a�:��޲�z\�.�Hx1�����r�m����W�]��C{�O7P'�t��'������3&FNYɛ�((Ĭ���>���◿�\r~Om��}s)E�o� �<�N�1���+��Ga�
C#04o�(LռJ�^��8a�8��!y��*Ͻi���1]�B����Ć�ͨ��`/��^{<��J>�P�eeĢ�_��y��s�8[�������	bfN9���햮&>
o~/'�����=�R\4��L�!�#���=�F�Ў �CY@��`vi0�2�|������V�R^�J�
짟~��՛��lP������nG{�#���2诧����_lz-M��7m�|���Y:#'���	��g�2.wJ_�U2��Yy*�~
^�a<��y�����GB7Ѿz��eedV�e:t��������U+ �Y���8�����U�KE��_��f:,DzH'���Xu-�i�4�J#0o���������3�k��Ϩ>����4�]��h����O?�-�6��C���c��)�����z���D�NV�R2쯺�*+���?h�b� ����}R<f�7o�;5~��Z\�P����8�#0P���7
�*������pԘ��
ho߃��_���/�9�$4�c��4u
N�>�N�2X���F&�c��{v��;��U�b����>_|!�?���GG�.lټ+W,C���+״�]��/��a��=hj��_��r�.��S*��6"�<�<I�JA@:���;����Yu$�>��
)�W��C�d���f�J��ߦ����o����ys�	�T��=���d��*b|�ᇍ+I-���,���=�C�,V���z\'������L��p(�DW�v�1i�4�{�\�&�F���� 	#��b��f'����y�e�+��6K�[�p��cxk3�a/�#G�!ѵ;wnF"�i���c��{W'��rؾ'���0>Jb6V�_�B�yK���ok���3 i�#�7}�C�."c%3�xi�io�3�t:C��#vx�W���2�L��� ���q�����yZ���v�a�
;�>NN+z��n�_���N��X�a!��g�KN6�ö�q$ytv�p���4������� V?��R:iI^�7�������s�W�y    IDATq��{�����
�|�tn���s�I�6)������=�شq;
�0�m�c�)s���Et���R N�.R�ra0����[p�h��j����xQD��t�!���n�7�Շ���5+^��N�\�l\3��#ͺ��ץ�;*rO�Y�7��Q9���?���[:gW�<���3��uQ�X�"
�����](ॗס��	�mÉ�N�o�d�ܼu�%�l۲���{�J.�\sK�����m��o������!��z�أ�~���nj[���g�9�|7�n_�L*iڸ?@n�6�����6�cܸ�֞Q��_���)[L�z�[�b@O���"sz��E�����:(�;yq���(��\��o�i����5��`P6�ܲT����O>e��dOe"��(���iՋ?�$}TIHw�S�ߋ���ں6mZ��nrd�ΐD2��ϯB0P�ݻ��|���~�2|�E?��f�Y���D^E���������f{{���}�l�Q��cƖ��W��p�ٳ�Iw`���Hg%��:;��~�&�|�X�������C�`o�(jt��[]T�Ϲe���i���L���RJ�����������P(�����P=�`��hY�1N\<ܣl���6�ai��ʑ���I��fNl]��Mvu�����˟��܃N����jlܸ�{��J��o+WmD6�Ggg;v����/C�%�o��k�������#�Jc��1����4��R�N�~��p֜���Ѷq5�.͓����q�m؂L&�u�:p�)g�{��y���;��'�D3��6w����L�`�L��9*4Sw�����{���{��4������¡r���_��/��]~�=Nk�,����~���]�� ��><f��x|�]�4i4ZZ�a��W�˧��`c�4��+���Ua���5���n�����;�������imn���n�y����������-�i>��`dK3��<^� F�jB�Ѝ�{�!���y}~?��3ؾmv�N`��$\�vK�$�3��\4�.�"q���ӭC�9�	�����;	�n��~�LM>���c��^�(��}�ڱQ��.��7~�������;�q�W�ޥb���g�q����E�̚�`i�3`���]X��"�TPc�捌��G���;;�ص�\x	�=�D�bx��p�-�X:���+e�Z��/ۇk��<A6
a޼K,�3�Ma�m��ٻ{��B��k��<�gG�6lC8ڈ��q�;'��o�TOQ=|�k_3�gF�z2ݓ�AGaB���~`1 /{���6���A�zd�܇�y�ߐ� ,�_���"�̦3�\bꕀPU.��ty��M7�d�B�5l۲{vmEGG;�9�����l�p��֬݀t*�+���ǌ����nK!��������o�����?P�o��#�3a�x��w!	��&���������Ĉ������Z1�ē���	��g������ގ���:�������N�nQ{V������K�ސU���uoٹ����j@��U�C�痦"�h/Į��^'KJǊ�[)�bB��\����MT0���(�v��y������y}��N[��Z�I[Ԇ��[���?�2AҎ�W�H(��TO+D�5��i�0F���K�E(��3a
O�/�@L����;��{Cc�&6�{;�ʚ�R�����uEE�)�j�#�@֬�-���zy8��_����g�{S{ϻ�1��w�m��T\T��I��S3"V�~���<��/�͛6��/����ծ�u*�A8�$S̘q2�u����mہ��zK3�{�R����y��?���R�7��ۀs���ݍk��N\tх��E0�����F�����{�PX���b�'a��3W����R5YuG��6	]=��ԧ,��_�2��f�i�`ж��|Ŭ��������ڜ��`�^���q1�	U`L�`p�L��t}��4����м.c*e8H#���ܔ]t\3���@J B�,��+}O�ϟJ���Ϟ=��*�CA}�(K���^>�hx{[r��#�c����	�us��GY�p��[Q>��_i���t�h<ԉ�?���ΝkkQ���i}�ƍ��̵*^)i�<O���֐�U�\o-���i��IF6Ї�s�g��SO-�K՜j\U��yb�<��wT��~��`��E�G�/�������'5s�?���bʔ)`;L�'A�}�9�=ʣ�c�����D�f�j���{�j�
[�&p�>���KQ_7d#(|����Z��b��c�����h�hR6g)V�lʢ�'N�n�܈�H��,��0�� ��"",��Հs۶mX�x�i��(h+ �����җ�d������Y���H���j=��{��*Ս ��w�۞�@��'P��gg��-p<�
��g�8Â�
��$�%W��o��o6�2��o�G$�]w�mD�e��w�	�����a��s$�x�)���i�eG3��T�Y)ܴ|Ư��e롯���~̸��n�^��nu�i~>�����M���c�# w�R$�2��*�'����-�%�sK�X�I�����2��J�*�4Shm{�y9�V����&��@��~�T 4�R~x-u�b^�O<a>u�[i��`�`�x��kM��t�R�df�=�̳x��l���
�����[��_��_mdAr<�'��'L��"�t⬝R��'.f���/��K+�;�S(�����/�ws<�q}%�_Ҝ�C!ׄ��/���/�	<j�X+��ĤS�=��ng�Z�Ҹz�z�ro�>���M���}C��Y=�<�pT��i��]o��4�ú���4<��;��P�������*�Z
L��XȦM���8�K����c��/8.�P�|�[߲":�6��κ�����y��n���sx��|�,
�����YL,ܡ�ƹ�Vʟ�'���P�'����:Ӧ5!W�c�����'>�ѣ� ݝt�鴍g>Wj���~�,zx12� ��"��&���4�\c}��$׮_��~�����3�
	�a�?�S����Ϳ��q�1��nPo�y_뀱�5ZT�����߼�M�b�}T����*;�DkF��K�Fp_�z��w�'�t*z,� `��:�ݏϨ����;�-�<y2����@��2�@��d&��h���x�������y���*��d�m�w���?�wį���<�M��/���b	���aĈQ&�#W��c�m�b�H\\�r���2k�,�`����	&4��{���{����a ���X��k��|j!��%���9K}-��	[�)]e%u��i����oV��y�j�/^���{���J_ڧ�Ҕ)|9����%
�4�e�!����q�Hx	�5��X 3�.����b4�K^��||^��8j��}w/��9�т��z;Ə��ꪘi�Ŝ�1A�߬�l��N��~�%K���b96����80퐂����y]�?߉���_X�̲�<<_��֯\�\���ϟ���>�ƕ��j>��y���J»�:��B�2d8��I(��k�YY@�5 k�d�RYܡ��^UV�u׾����rl���%v����*� ���SӦ��jL�:3N�i����Z�\�(�
ؽ{�Y�_|˖/�`�Yxp��IH�ߧX,f�[Zo���^6�����W�` l����h;%-?2���}���b�č� 087�|y\�
Ԋ�� C�+]�r��Փ��:s�L+�b�@n-�}�C=4K���"?�Lpj`|~� ��ǟ\���h�`z%�g������ K��UV�5k
��AG�$�;��I��97��xg�mJ����^ם�W�����1�t������T\O�J��}!�PЇ�G�D,Ze׬��3��s���Z�w2�l=���� 	���"1#���lr����u(5>r7�
'6$Rq��Fg/�*�D����1�y�ǖ ���WZyA��N��8����\^|^^��*/[��x���Z��ť�����.Ɯ9s��X������~r�0�DE���U# ˓���pMM-fgry
��)���q�;�]��/ 
�?�p�T_�Kk�����{��_d�h���v6n�w��:l��6`�~̂�a�	|4u��5�F޹���h\,��c0�~UnP��e��dpL����IVgi[�78d�3���M��Lݔ����H3���+�?e-�R��@����~�^KMA`>���	�y�,+l���u��y׊e����r!�{�����5�.���u�}|��<�"Zʱs�Nz|���[��Cw:�T&mY�W�;m��#����!!dq-�)�l�("UQ*~'A�FD;�#���Z�^7��-ŀ�:Ї�?݈��y��'��\^��)6����-�,^�1�Ә�8a�Cʅ�C9�P�"�����82�ɖ�,�8]|ʝ����&L�0wkIY�4�C�_I�/2G��l	���}6�����28_A �w� ~�}9�o�<��XNjE�C�'5f|����P������O��@��p}/_����ƔF#w��@��m�k�C��8�jb�ո�	�x/�W���'���=�Q�,�L��|yms[T����+뽏6�4P��xm���_
Z(���x�Q�o?y}9㓊R������w3Ѐ�(|�XЕL"�ݍ��%BB>�57|F>��G�{��=��Wf�U��?�nP�}Ya��������;�0J���T�Lk��O�TP_{�{}	cY\����|?zo)�^+���|q�r��w���|���:�ڰ���,Θ���w�Wpk���ܰ�C�8>-�XUM)�9�B�Y���ks�u����@n��>���Uޏ_q%߾>��O����j>.�o~�.�\^��b�t�wmmm��HM�	�|z�q�ۥ�b����w>������c�F���8&qӊ�n|����&PB�2���9����
��	��1�j�����	_�ц�������]6P_�� �E#`?	�;ݎ��,A�� ��է2�}��V�[��|pL-1@<��2�4~���ZEWy�5�׼{�Mq�}
��ރ�Y�W�e-����y���t��Zpoփ�8�R�O��SƞR_��y�A���[0�g�xǵ�|�}�������k�k���11��c��w �G�r��R��w����'�&��f���iԇ�k���m����*ȕ4z�p��#����������Q;��W�ل�G �{�B	�$ zP��i7�_6�����{+��9���WC�����aN��{�B���L!fŰBPy��'�Ng|mK�������b�U��S�0���@�����;�C��k����iT����*��c=އ!Ϳ�ٚ�`�/�����^�/W�4x�b�?X
ZQ�C�!�]�J���K�0y}d�݆����}�f=�s�ұ\��E2�EE��"X6Iݜ���S^�}	�y]� �==ǻ�D>�5��o<�~Me��_�����p�L���h{�Y���8��K�;�w�Cm^��R�@~�ײ��!�?����>N���t���b)�3�C� ���>�`	&�B5����|�S!69���A�?�~_�P�˗�*X�0�$ �R�	�S�2�5��e_4����!�?|��/*��}z�?��l���3�K�O#������p.������e�x����W
��J@����A��3o@Ϳ�p9��.�n�G� C����uL_i}"�� P���ؕ�/����^�UX�C����:ʜ�ޚ����3��f���r�i�o�n9�{[O<z>����{�!�<���_(��1��7����qzh�;I�$	 �M)�._7d.Vs*7��+����a��}\@]�CK����+�?}��Z:�?h�>ݩ��;P�t�!�?p�}�a½�z����U1�� ��-����[���om��`��-X���x��*���A��9_�:���W1o��0&�������h
�L.�M��������G#~�@��+Ư"Q7�U���U,���7j(e�0E���������"P�~��������ZB���R�?��q�|t�Z<��*�Qі\i,2�Y6W��Ze����y.�->�ݔ���1�G�����0�^�z-C�S E�9s�(�O�U9����nx�p�d7�錍m&�~P	QV�����|V�6���J�9Q"��p��*k��s<ʬ��b�bU^
�ǎ���X�� �k<�TZSz{+�5��ޞ���Y�益=�{C�Z�'�jo�^Q���G�\�-aV\>_N�渲��\=~ �h����=v�+N̻b�e˞7�qWp6��?��y�"���������q�?W��E.m?F�����zm���>V�=�B!���&-�j`�&K��k�8��*�i���#��?��% T0t8��\�L	�ci���w������n,��R+T��Whv�L�6���U9����K'皙x+O�!is�oW8�tm`iS(�"/���=^��J�������E�+$^���������r�����@��)巪^�hir�Q�H��.9��8q���lh̩�X�TI��
�%�����sz]���~����|g��8�t�QPp���sq�xoS�I��kk]��������)o�s/�'��Ϥ�=�i�ڐ��U��.\GV�۝Fsc�1�2|ذ$Sd�u䆉�k��V�$�[���9\�\M<�p���/��m,G�Jt9���g�y.�{>��r�O:�4nFiuiv_�۷�4C
m i*� "��F!�	���w/�x�B�`��F"�i�RW�~��/�1I�Tۻ��	��	V��x��}P���N�J�7 ���#F�w��W��ss.�R)mb�8���;����x
x�Yc-�d667�S��ל���_ȣ:Ve�.���pu �Q4��
"�c���Y.���������:3-��E�,&	6�#��(���	N	X�{�ݏs�{h�Er�k�;����Ha�߇�E��,-	j��Ƿ��ގ�=^
/��'��s%���g���0�Z���ӊ>aډ�����W�.�h4�ؾ�:s���T�zV�X���q�Q��-�@�ɞ���/����x��>�>$v�3kcU��e�I3��oKS#2���X��Yk�F�-.��ԩS1i���k���.l�B�a.|.n�#�<�ƍ3ӍVB���M$-�C�?�:��~ ��MWGg���h��_<�V�	ۻ����{r3�1������ �U�oV��m�L1	g��ZB��TE@o�W�KSK�Ϳ�CZ��xe�\�Qy���w|G�]���Z���ޝ�_Ȥ��҄=#���]���=w����!��RG����f-!���Xr\ml
���:+a*ˇ���J�)	yZd^b;���8n|w�I�=	��LyǕ�	]�	bY�K�P�{o�Y�)���:֫��~N�:�����~�s����r��9%(�F���q�U{đ�DB�fRض};�y�i�w��Z�Ţ��;|�H{�h�Ŀ�?��'k�h�i n�A����a<�qc�oմ����q��ދ�G����(���c�`˖Mf��������Gy��v2b���nH�L�~�7qQ���<�_c�@n"i�2����5�v�����˟1o�E��H���|�I<��2[%��ߩu^xᅶ���
8R+	@���&�Q�)���x��)�i���8q�]OZ�W�P�}�=�II���^b.�#�l�C�^j���e��r�xP�����;y�P��B-͍��c�8��+7倾�]1�<y�]w݅�/�����F&H��ƙk��#8_����[��yK_x�>�h��D+�q�e��36GlIK^S�7ޗ�p�w�y�)Di�_��O9���J4^��uE�C6���l�Ə,$�}8FrG��ټEc��,Y�[n��L�,�X<F���1a�8�
i��	,~)^Y���&0�!\g��L���3g[G&<��_����j��F^\�7�s���?h��?�'�S�.����w酸���+f�N%�f��xa��,(GL�O-lW{J��s    IDAT��������r�����F�L'����6�}�Y�[��� �!7�c�=f���J�����;�k{�K�5Ea�9�6��K�$���{���\m�����5�\c��X�x�cC3�{��6m�\�*�F�v+-��8y�d�i�r+�Y�.
�qd�1���K�N�/�7�bw,cW,���s����c�<�쬪��N���IH!	%4�]P��2"��"
D�*���S��\D)6H �t, ��i�L&m2s��~������̙3%���'�̜����~������Q���ި a��}6��{�=���FΪ�j�p�~����4Z>��#�;�����f���Bs�8���2^��/Y�T[.ug��Y�|G�\g�64���˵��|3~uS��ڧ��ֲ�Ro��#���4S�Y����9R��q{)��T�E<�|����i�(Bt�y;J��J>�!y�'���u��qo(�\p��Cy�S��?����V��{
��"�3�.���mr��G��%y��X��t��Z	8���e$��� �l�Pe�w�o&��^q��2k��2]��c�� i@���Δ��6Y�r��tw���<��w&,�ΐ�9�<6��p�X�[@�Əf��~�i�%Lb����!|m�r�є�i�����y�W�blsr���qPbl�{u_ɺ1��5`��f7���D�E	��ۢ+��h�ԼV��i��9�����g��5��� �W~�����C�h۠F{�6|(���i9h� �O`�`lX�?��������t���K/��ӧ�����k�W� *��oֱ�/���	L���s�Ygi�l���1�e�*T��9��́�N�lNۏ�X9�kZ��0��DkHU���|�u�i���|��k�T�� �Fu۫~�k�g�ش{�=���|E׽�]�y��=~?��hw{>�=~�}③ll^,�T�������˜#�X�(/��5M�$���u媫>&3g�.�lA�x�or�=�H,��}n};#]��~[2��J�j�O�� ���ڨ�}�r�����r�rI��f-�M�NGd��9��cK}h�������	�S����Р��CM��S���3��r�����8E��̵r���1c�>����#o�q��hO �i{h~F�������K��u�P7���q�  |��6W�k��J1�b�?�^54f�Q������yJ4E��q��&(��Z�v���_j�E����瞳w�/�P��t����E8��Tł������ G�q^�*��;�MPs ���35�ߴ}s�+�Qp�6��)SJ��	_w�y�j��h��Dw���t6�6׀?=|�^0��7ø�m��+��_���9��W���UysچR���i���ӟ�eie�yN�w��Hn�g�zHƍ�˸	�d����U��tN�-]-�\X:�S�����sϒQc��ˋ^����_��͙;��ɶ�+�?�3,�ٻ�&W_�!���ic�<���r�GK>�%MkWIgW�ĢԨ��斤4�k�l6&���d���Ҳ����җ���'�E�hٴ,$۴��'NP�0-�4EӺ�Kܞ��s����cƨ�vb �wM�t�E��pԨ�ȖIH�ײV���h�f�"�\ )���`416\_Z�?�/�B�'�d=�����E��s~��|l�an�]��/��8-LШjh �1�t���CF��o�k��8�]��q2f�o�ͥY<G��9}���ic�o��8KN�~�X���J�w��-��x�W��u{��W��c���uO�ߡ�� ;��{��gk羦&GU�u��O|B��|�+�'#���3F�,}��ڰ'��c����"�iiMI,Q/����$D�I.�ma0{��l���G��?g��&����G��s���#WX"�����By�O�!��-�XA֬]�m1�
��l��.�6�O�F^^�V=�(�B�(,P8bQ$��pL�����Xx�Y4A5����4__s5A��-n�O7��1�	Rv^�����67	b�e���>��kn}�ôG]��xWz�:��1���� b�c�����>����S>���'��ρ%,q�\�:��U>��/�?��aB����� >���O�z�{3Kz{��Ӭu��>�\N#�h�������{�.8}�~��l}A�]q�J�-_��<��{�G�'Ə����)Ţ�ĥ�+/˗5)�l��)�Z;��o�Pԅ��䎟Ȋe�J}�s[�����j�Oz5u�NS��k>.�b^��.��m��c�L�]6nZ+�=�.����d�4��$�y�ؒ��{�E���*~4>�i4`�J�^8M8P�p���;��1���Ȩ��6y{.�j�f��Z�@�`*�8L�y��}��7�EE��iަ���>3���=�����;����Aɿ�	=�,�����ܒ���(�&����k�v.��]���+ 6���o�3��M �
�	�Jc���߿��*�����s�������2����� ������Ϗh(�2���X�PfX(��׭�'{P޲�,i�8ZV�y]2� ?#��lFd�+�K$Z/�YIeC��]'��Uo��fY�b����R�Ap�������i��}��1r��?*�u52nL�,��Sy�>�J����u���ۥ�G�	i� �[��+#k�&��S標�Åޙ?~ɁH��SN9E��Ǎ�R��[nѰP��\t�F[����j��&f,o4�������L0��i���f��`?_�5'���K�F<�}4��9���h����(�Uic��H����l�|6�v�6�c�='��} �4�V�Uc��߿����)��l��������}'�/��y�fY�M���j�f�� ����9��w,,z_��X|��ΎM��ӏ�N�GI"�ի_�Tڕ�A{OO^^|a�D�d���r�ۏ�y��֤?��w/���������3�gvĂ�i�7~��-yU%ڇ�Y��Qrּyr�[����VI&7�����"�0 �➡~��Y׼Q�6o�T:$W|�*}`<�[o�U����׿��=1�h�\r���%�m���.�C��k	_��,zc�x8�/�\��4/_����/[���[>0�Z5�� ��7 �/��|喏��]������<>�җUe��K8�}k������J��ӷ<�}_Y�����6��/��p�z��Z�׵G~��7_�~"��?�|����͊�Ә��@���j����ѾQ2�N��R��C�����BL򹰼��5iK���^";�<SCA~�a���%��T��w��u�=w�}{����/���xC�=ye%�ϓ��T�n��v�X$������MR�Nm���K!�x�N�;�p�m�=�D7�勉ǂ��K������w����%���A9j��x㍚d�S_���y0���Q9�].��V3�r-��r@,�0 ���%`/&tʩ!Ӽ����W�����������2��}��\�3��e�F9��[ff��c����W����TK4�ݗou���r_�9�4}�����$`����Ja��l��K�'���p?����K.��2I��*���חȚ����t9k�#TN$��ttfd�Y��A���@$:.��^eFՎ���77�a�e��Ͽmā�$/�_#k�9�t֙g�	�'�I��Eem�Jy��G�E�4��E���C<DN8�d�0q���&����s>��'1���Q��	���-Ġ_w�u�v]�j˖-�gc��e��+4��6������26g_Ԑi���� �\s���G����1����s�F]�w}�5|����[�3��)��@����?._A(�r��`�mǚ 1N��90������1�[}��h?b�W ����XC�w�;\ߊ��Ӭs�s���WK�K�dlD�� ��<���}�{�+�|��c��j��_�����4�]��� ��g��M�9��s�}$�/j��G{T��կt�`�/pM����M��p����dā�����f���*���k�/��޲�d�i�0�����.kׯ�H$�^���Q�'���x�F�v{�-�76 ��,��,:�a4��{�q�>,6?m~��w�߷LO�2��6�m�j������V�7ЄmL�¡ڵ�|>�����7�-_p�S��P�Y۹lN�D2~8����1�9-⬿5�h�Z���i���ߟ�r���{���)�}�A���5���kв����w��cʬL���a��E5���:���.3w�x$*�|J�I(]�\-�J��<C����Db���勲x�k��L:���Ek)���;�~������)h	�?$17gyW���c�	z�n3R,��ڶ�X��H\6lؤ�(�`8{��q�<c
�>?1�"�.]*].�Ӿc��@o8����w�\����\��U��>ܱ�����w���	Z��\)�u[i>�\>������KHM8p.~�4q��}�9��{Hm]��pF�Ơ�s���W���ߟ����w�a�}/����
`���T؍	r�TzB�ϸ����d�ӴD ��<$.��W˚5k4-�� �Gc8�st!|�ߔw��r�W��C�_��7!�?����0��l���\~��-^~�9c��(�.�n�3���1��3P�ӱX |ƌ�g�$.�x�����߯`mt��[��:;z�V>��#d֮��J��m<�%�)����/��ؼ~�
����:�{�
��Xο��kRa�]c�b�uM@��3g�t��ٔ
2��E ��n�KI7��'�"c��D�|�T���p��iZ������V��b|4���YMPq�JiB���m5���1�n3`����ӸSj�S����Z�T�%�+�}OUU�^@�6|��h9�F���)Sd�3�&Ӓdv�x}�J� l�����ߜ���\�ol�)ٞ��R��{(��n�� ЇM���+�f�?U+�j�HfK�e�=��h��=���t ,�`���{�Z��~D~��ȢE�Jac`���l�d5�,�6����T���lc�{ ��ߎ�7��~f�PoW"���ֱ�O=�TU��A�ɜ��`��?�h��|�8w-��)���}��8��	ܾS�x9��jUϑ��6sa.�9����s�Ľ{ci�����a��s�2~��7��Q>�yv�Z�.b�����'�"ف<d���z�qu���ʬs��E�7i\���6�q��ގ�w�j��MX0C���Z�r������O�'�?��u3�9W�y�1\3 ^vL$���G��� ���w�+�F��?w���d���4<��SIO�>�$�o�]X[X ��kSP���9UM�дa���Z�2�V��pJ>x�AB"Na�},���!}����i�&��~�-.,�-��������������3��g_X2�%l�!��\����J)=y���{���U�H6�@�I8fmb�*KmM�*\q�Ǚ�^��M;�#B��#����xK�=yI%��|>� O{�z�Eh◭T��{�("�|o-u����� ��_ViM���a�QŐ���'�/�o�m�X��p��%�X}|?���E2X�J���p���;f��},`¢x�ꯖ=nܻM��('����5�q���Vp>�f:�v�D��������Wp/��\��B���,��3�4�������8�*�O�n,��F D� ~H�0���F�
���j�Y�u�c��'�.�����c�@����]�\��Ec��p7����#�4ݓ�s�Q?�EE(p,��M��Ꭳ��{�՜&D���1#��}y�m��a�zO)ʡ �bX����tc�z<7֓����	u��w���T�����g�r%,"N�{�iڼ i��^�Z�
7
��7�Is��G��d�?tE���\�4��
��.�;�R��Pi&�����c
"L�N2 ⺨9M\�GhX�
 ^V����
)dz%�����m�2�/+�ZB�{�k����Z�6���4�+>t����Pi)���L^���9��SUU_4�5Kry�21*E���D����x4��H��Hb���9��3���MH�<�Ũz���ϲ��֞�H��	�hB�Ǣa����ϥ�~�K졭g��o�˜�VEV�� yʀ�֥�_�)��o���xn�G�>2���
Ղ2S�d�}��P>4��!3�%�0.	���}O�\�v��sP�G6�W��#!��b��$1�,�6��� �Y�]X�E��D
���F�����-��s���?f�I'�K�w�y������ӱ�5	m��|J��X �>������n2�`&��8Z2y���$�1	�3�tHM�[:�֋d���HݨIR��%��c"9"������ϰ�Q	SS�%ߛ���l�N
Q�LT�y�Q+�ܲ^6nZ��^5-�C���~��d�`��VdN�.�ϱ+�3�����7!�X,��>��-�ʔ9W&ȸ�j���;����p��l�Y��`���9����0]��J�*�|���?�aҥ#��Ϗڒ��*i�L:@��C����a�e2���������g6�.Y�����r��6�Z�v�g�;K�O+8�
y��@�i��o���f��_��u����/
�c)�$ �m� u6��SN9I�<{���Qb##�IL2�uHw�
y��dݚ5���mǾSƌ�(�bA�E<�0�XC �<�
��Diբt��k$'��8I�k$��H1&ɶ6y�OԒ݉�:�Td���/p��̙��YT�$�Ȣ�,�k����O�����DùJ��	'����{�Z.e�s�b��}�����e>=��h��M(���zA�%��{4H�T+.PB��2A����_-��'~�i���k�FMM�F�(؇c[4Y/E�� �B�F���˼���n���P�M�I�Nш��e`<�̢��;��=)��Iy��h�#l��\;�l��Xb���!���*�l��J�G
R�I$�*��:���Ț�Kd����ݍg�����y���6�m��d�*Z�)���J6:^�?C�z���i�I�������vB��'�r�c�� @ȳ:�3�$	�>t�	&@��}[so���$f�(�ǀ�$
�q��aaS�B��������؀0N^��P= /�5��C�R?fQ���2�SJ�?��[]�o�4��YҹZUOʹ�)�ȡ���ۅ[9n������b��L������+�V�i�,Q*%�˨��F]�Z ��S)�ɤU��L�H���t���-5��&"�#t(
Ю	����{�±Z܊��D� �\���I"�"�^p�lްF� O>�Q����G�F���ry=����c�}$"�P��#�$/����-H}�hy�EjE�ui�x�s��{�� {Y�y��2�47'�>3���g�f ��Y�Ͼ�i�n��O"��XY��7�կ�ϱ��@ྍRV��r�Vp�ņr��ou����J#	8��ܵ���c����;��dۇ*�>,>�4��:�ҮA3�#�6���w�}4������
h"h&hZ<L4��1���M|���|�v��U���%�؈�	G$_�jr�Y/�x��82���wu���qN`C�`��c�f=|�J���*d�.���P��:W�}w�"��keڔ�2g��R;a���Tt�`�/�׹�)�~V�DX#��IE�J66Vr����b�F��H��I:�s�x�|U��P�7��8�h�Dv�\Y�4�ӟ������cL�5���&�:�,�����k������?�W�u8���-�����d���RS�ڻ����h�
���~�D\B&�SkE��׈�j�����N4�|XT�pL::�d��3��w��͘Q���1Rp��ާ�|w�,>�i4�%����Oߏ@���Q*��%w�_�K,'s&eD�D��gs8<��Y%C;@�0�H���p����3��)��&��i�f;%�k�����n���52i�$y׻eB�N��I�)��I<�W�@�O\�֑��|1,�P\ґ1��-    IDAT����Lx�d���
jRc��7|O��Z�B��r,�2��G{Qd2
 &<�֦�����G}���e�����G�{${�,n��u�ܹ��'��)K�B�ׯ�iJ�P�����Q=%� ��!��|��r�1����SU1����ē�* ��]J��T{�#��5p'�V�,׏�M���#o{�12��4M��f{4�C��_A('��P(��1��'�����vg��o�|���a����z��|Njh�I�i��pF�|�'`�!�i$'E�hS�lЧ ��n����@ ����,�^�7~�g��F!-�BJŤHO��������2m�t9餹�0e�tt[xja����POH�BB��h�9�	�M�j$����z�>C�߰a��薛�E/�0@�V�۞ c9! �瞫�}ӊx�-&h�ϛ��|� (�ƽX3h
�)��Q�*f{=#��L�(:m��ɹ眧U=�����&�F՗rn ����0�A::����ğ�T����j�/��dD�>��������G+�>x���h������|@b���]'==���+�i�Ji�h�D̳=��Kf�ds$m�f�7�t�.V���o}?���4����[5I�c~=�<��-�J��R���-?Q�?����Ȼ�}ݜ ~�����$���4�����w{�?��X]7��#��vi�u-ᨙ.��%^h�pz�ܿ��Ҳ�I�N�*'�|�����d�]D$L@��7�gP?�����? �/D%��tt�d��[/�P�&|��ٞ��������R�\���@��̔+��s���a�DЖO9�Ufx�[���<s�G��5i�ja�>�VC������k�[	��4t:pN�x��ަ�N3���e���I��J(pN�)@�˚�����YH�ͭ��ZP���=r,����#{��C-r�N�;Zeٲ%���0y��m�=eԘ��Jgg(�L��ؔG�Z.�F4��il�v�=��J����l&/ӧN���u���mw3v��\�T^~�yy�����E�A�%@gƴ�e�}���;Z(���z��'���]�t��g��P<���L^� <m��kl����a��5�7Ż��U	�K����$�RISP�����XM��p��%W�v���I1�)5�#��&��*���Ҳa�����O��:�cͻ0ϡ�4r)� ��>�� Ӝ�I&2�9|#��KǶX,!=]���?��!I�9�a8�>>�E��U�X8"d�J$�O���0��#�=��$�
eb˾cc亥���w;�ʐ�&K�4(,�p�PO4� }�#?��?��pn���_�Ĭ{�@Y�2������n�:�h��y���?��J;�C5�1�M��e��瞑�uM�A��tugd�]f�G-�춇��.��GV�m���9��w�?����B#jf��lZ
��,ym���ҳR(f�.�~�$�HWGJ:;3�����G��
��w��]u�(؄���g��?��j.<0u�i������g�yF��玚��x���P���L$H�l������m������s��(��P�S��Pf���[�e�j����j�)�?�揀��Z�B��֬Dk�P�JN�%������	��p�v�wȝ?��<�ğ�TW����۠% ����I�����wb�)*� D��c�t_����+Y`
ʶ�~�������������}�$Q��c��|���dJA�B�/0�J1�W'k&S����䢋��C�=�~g�)�����ַt�~tc����_�4l�����^��^]$�m%�^'��:I�����#�~�z��݋P��]?W_ k����0i�#2�s��9�J&�?^I�g�y_{����.�fH,"����"�F'��e��l^/==��$��rE�ܒ��%3r��)S�(x[M��i
\�f�Gu�nD��X��K��అl�}�-��K�`J����$�$ �A�
��)���}
P��JZl/��UMG���4v��%����������e'h�������0��|�o!\�"Ų$_�s�ђz�6qٸ~��z�O��?�4�m��e c`n`=����k����g�r�Ъ�<+V�(Պ1+´c�?h�"4��-4gֿi�f���l��QF	��Ϛ5���D׻��V>�����Y�k�>X����(c�D0�P�$��{�{�k_�����8���.�HA���p��4��/�X9�I�tHrs���6˺uM
�(A�C�>���^�^:���K�a�Nz����k�#�}�'ߑ�z���%���l~^�N����5��6�{���v���e��W��#��_$��u�7K�ڍR��,[�^�9��ڸ�M�"�����d�����f8���|�C�/}�K��iM)k�q�8���CY��!��d���z-E��8οv��
��2�k���u�����餝�{�	�L;%Z�,��*���M��NS�?N�'c'L�t7��f���߬\��a�0GaM��b.�%%��d���ʈD��i���G?�%˖J��m�/�P�`�_�������X)�A�Y_����΍ՊF9m�4}ˀj��9�ǚ��?������6 h��Y066�T�S&�	]�N�6V�p^&P̪�s��u�]'+�-�4�cY��%���|�;
�P@|n>����o!-}��2u�x�PN^}�F���¡���s��2v�N�t�j9�'ɻO��x�Ң�jo�,ݻ��_O;���/�s3��,���c"��l��$���r���b�G6�4K{{��c%.�iY�n��sY��]v�uO�n?��M��/|��ݢ�������8�8|>�я
-�xX��o�߰�]�~�W<�ޠ������Z �_5�=�/�w����U6KK���c]���'�3�����e�r�#�|U�'��������t�<3q��)��eu��3;Dy��D]M]��Ʉj�G�K6<J2E���g�f�*��?��Mͮ�S�(7��_�y}[�?y&֏��8��;�	 �~XVn[�&\��� 5����8�aj~��9�� ��bV�YF��=7� �?zf��뚀5*�_��<��g�^��Nj,z�(=�Qj�~�U�Ę�@��n^/O>z���,;�N���AW�?&ٌ��Eˤ�v�4��$u���ǯ�V��FIgw�^kŊ�zn~�����h�l�0�k���CW^!�pQV�\*?�k9��äP��VKWW�s��jd��ViZ�IB�zY�z���!�)g&�5�\SZ�,z{8ַ�
��ޟ$R��8�m�9}�`���s>��� V����5�	p�u���o��匇�EI��֑���
:�!
B-f$�k�Da��3����&�}��ɪ�O�?$!AcZ�?�H�\J���7,�bL���;!���_�1 v��%Z�aS[�UE%t����mƀ&b/Ӝ�Й��|�R�P�7��zt������$8z˜�s����\�	�q� �����H;�()s��}[�:�F�"�L�.9�i�t��gȧ>�)u�ҫ��k�U`��K�B��&�h�x��e��k/���J�<r_i�4V����1���l떥˚%-׷KgwV��m�caٴ�EE�.ݲ_���Vf�h(4�=gϖ�\}�Ĵ�C�����;�y���]�~�jimkQ隈�K��NY�z��r1y}M��e߃T�ǼE�n�Q�>X��ӊS���Ik(���g	/��@7�v�cK�qmAT?����\2W��?�}�� JNi����^�+ڡC�������?�q�u��LN<��D�K������|�.��?~��h4RD"�!j�Nϗ��d%$4 ������}����#	��(1��|G�l��5Do�������M��F� �ti@���}�!��1^>?�uW~,�e�o�I����_�m��˵�"0G��6?�o%�IO��í�i�Ҵ}_0r?8|���<��#�<R-�;�C�.]�S��g�(�����<����̖q�G�kK��K��D��saye�r���ٕ�L6,���:=j�tv���C��0&?:�����n���5�5������~L�j*f����ˡ�'�b��Z�B
���i��M����뫤�#/k��ȱǟ��?���8�j4R1G�q�<,6+&�]w�UJ��}����M��^��m?k:R�R�4.��k`rSBAk�����x�C��崺'��2�
�E��ˠ����Z��K��#WKD���f%�k�p�E��M�o��u�d��i��O��JW� ��GjS�;res���Y<9��\l���%-=��C5�'��W_����/k}�����WU��d���b�ͱ�),�}_\������[Pۦ���%
ڒ�ݞ/�K@���S��,��^������Fa��^��P�,��PV���8� �gs�Z����(k��a��iz]:�h�p8"�]=�|�jIeD6o�:\�8���+�_[.w-�/�5�m6���ܹ��L�]]���]�F�{�{������ukVJwOR�6��\�Gyr�$ź��U�o��Y���רs�ŀ���4v��v�J�{�WZ���A{D`��㎅R��s\s�j�O;.��JN Zd,���u�>���xc�����Ւ��q�:)3D�E���u�jA�l6%�t�$�Ih�g�Hj�<xϝҺa�L�� '��Q�O�.�T�GE����{�i���	z5��aL.2Z
�1Z�!-5"�z�<����_��������C���F�;��sh���r���A�<���a�>5����l�}��6����oK>M��K��l�K֭}U2=mZͶe�&���n�hm]��^�$[���ʵr��W�����p�N~��?�/�KF�%����m��8���m��+���ƙTJ�._���$P��d媥�|��QL*,�t��5������3%��V�1swV$?mq�qN�iF�C��x�%n�E�B�s˜J��ETqkT a�泙��:���db�5;1W�=�5�kj��'%�Z7��U��?�u~��-k��1�[�y��w ���F�eR��vK,��!�l����r��ۥ�y�4L/���4��O��H������<���2�4²q�a)(��B�^r�1*z
1	'F�g�)��w�-���Ev�?�����/�}i��Q@��?��X8u�@���9�9���/��ژ�3�����M��A	%�GK8�q���7ȸ���N)Ƥ�'#>�;��?�s��~��ɫJUϠ�b>���cG�YgΓ�;X�]�m��i���7JG[Ri�P!$�h\�L�*���Qv�6K+C"�)��׿�����x8�}48U� � ���4�����kU��*�O��q����Z0*��%�i�OKWG�߸�E����$	�Õd#;���@�/���S��f.��{�w��х|F����%%�L����_�*�Vj�ƹ�d���E���lZ�ZVZ�IT{���/��/���I12Jr�Z�)F%�-�L^�Q��ǷH"�V�v���b���,D��2F��GI�)�����w�h�믿^�=`N��7�B&5��x,,�L�<��S���OHw��E�g����Ւ��s̱�����3V��^�Q_KJ���������++i�tɱH���0I�s�<y�[���DL��Z6o�H��+V�����HmM��7^r���?�L���ø@�RY$h�˖-�Tp�r%j��vq왃W��ΰ��_� s�r��O>Y#���:"�Y�+�fZ|�UWT�z�5�O�1��<�v8���N�����*g�{��I!��P!-�ѼD�ݒ�l��~�lni��;M���q�$�FK���Dj���ϕF8�5��/Z<>�0��:)D�$NH�>��:���R����)��H��ڧ�2�w��ه~�nԜ�D�QR�`�|nV?�d��Ib�߽�ҋe��	l5��sҶy�,Z���\�R�'64(1z�X]�������=��qB>��_��?w����+*�?tN	�pxf���w�q���{�)��u����%� �ߵ�u��IgSZm�����-�>Rn-��+��� "p�P��/�+�A����í����ꩧ
U�Jt�g�����|�s��д,�?��I�=�y}���~*�%�&M��ft�m⡜�r)I�Ҳ�y�!p���S����K��ه��O5h��<��#T �HB��I���ȑmIm�M�em�j O���Ù�ߡ�7[o{p��c>9����M�+�y����^�����l��o�8�!� ��sl6�ў�T�em�_9.��+��������Sa��1�uw�q����46ޔlO^^	���IM����Ak�\CC�w�}�|��%��C(�鲓��K�_��,~���q�\�߉r �k�]w������H j��3����@�[4�j�A�ᆪq.�K��h��VD�B�}�1b���E�S�`�M�X9�� �j�ѨjN�\A{&S<-��Z^
�n���G�R[C7��� U"q���?Q���$��Ȃ���91�XH�X����G&�W�N)�"�R	�X�n��/�},J�֩	�сo��/L @�@����~s}�].��6N�i�2(��f�TAA�US����fy������N�����r��i���8����HX,��.$+���̓�8q��;Fv�4YƎ'�LQZ[��ҲY6on��x��f|FA�h���O>���illT��駟Bİ
 ( �~�����G/m`n�DS����@�NA��k]i�����s�nL���D#��N1��
��pQ��٣ɴh���ҔF����fc�*�e�xI�Y�G4Ɯ>�Ez�F�bk4^��c��3��(��ZKH��[�C��ܕs{i���\@ohhJ5`�*{��k�.�{([w�y���`_�P�~�����t�"�&V�J�n���"��YY�v��X�\�֮�J���Je8�S.���z'�[�gNc�-���%�4�^�ؚ��"�J@K@� +@`��"���ʩZh��l~��Ԇ�BVl�c�.���`IahF�{ktMY7��(����B���-�6���)�ઍ��E1��r���"EpÚ�[Q���h������x�P�P@e!����I|ύ��U*a�`�--����`q�V��O������'�Y��	|�����Lk-�vMS��������5�<[�4i?1��k�߯Y�ܧi�(Y�� ��Z�~�i����I�$w���to�M��?�>�����̿u]3!���YG+\�a���^T_#�g����Ȏ�N^CE��j�P��ҕ9��<@��tJ�o���n&Ο�Ë��;�s4������Jv��	zr�i�Gi����F� ��Z>����| �WH��m���!� %�+p/}��n��p^.z� 	������%V/ޢN|�|�1XL��s~9 ��FeP�pŅ ���=h$��mnݢ"��Kz,�B.�^B΄{�롅㿢�N�����˪�Z9
n5���z�)���u����_�@m�@f��,q�G�PG�:��h�֢p�X������2��:��]�����ޖ�����ی�i��)�
�1���p1@ӌ� �@���O'Q?<|8?٢p�֤�<�[h^��]��Uz ���瀻W�@_-�-^[&ܠǀ+��ZVV��IT�e-�$z_N������c����7��'�O�:a}�R��i���[-״{��
h�\ֵ�t����,b�Y��+_<�ׅ�|���z_`��û���,�J�P[�(W��qƫ 3kz��a1�~��&J�T�=|���A�?�A9�c��K/U@�o�x8A��"G�h�Czq��r0ƔI���}�`D��@i5�Kt�o�M;���(�JZ�3�\sj��X�l(8@�l67�  O��
�ق��P�[]4�7��0���5|[ݴ�ܒ�\��`ӻ�x	���m�KTSp�����?98�X7Dy����~&����5��E�JQ;[�oL)��>��iHBt�����n��Ÿ�H�p��j���:�4�H    IDAT^6�����2�+�5�K�'9�zDd��b��c�ҺY��j�X�{3��"�'d᳧���Ju�Z}.:���#��t�9x�G��6�6Wt��+; ��`�=[�}|�|;��_�K���7.��V`����n'��3Yՙ��d����fZ�{u�Z��>ڲU[��>�?X�zەuc�����7x'h���m�WI�!ʧwc��p��1�w[��J���T^Vc��%�k��_恵u�ŗh�M>���&	���
�Ma�3a@EJ4U�	pn�QiBd@�Fnf������)��oq/�X�:��t����S���1�����o�� 0��>y��'T`�z��h����"�����E�Q{<C+�`֎�OF��C�I/]��:sQy�·o�c�>[������ι9�l��o��  ���X���p �x����X,�.O?�^~��׭ҡ�c@0��g�}s���������ӁƯ1��a�Q��������"��G���;�('�P��pf������b@�o��
��'��¾l��Y�uiA�Cz����}�l ��?�x	p��d��p֟�S�'%��G������W��͌lo��Qg��4wb�*X 4�D�'���R���_�}�����@@���9��}� v@��G���ZtE��� �~���V� ���<��C=u�IL�s&�h�����O����eԉ/ }��Ea�ꄘ�"8,��L��/��m�;�;�T���
4P�Y̹:,:�D��:�0V;�؂�q�����cJ�O4`ͽ����;�*�"
(� �D����o�� �w`���h����?�.��q5˭��ӈ(p�B5RR���&�O82�o �y-'d8�i`��O�:���&*f��U}���n_����e��$�@���k�6�̀�5��B7�۲�}F@��7��+&<��nA�8G��=VYw�y�Sm���f.�&y��O����������MJ�b�3������a��LR�ke!�>�lQ[g�;�/�7���J����~| >�n�(e�z��Q5��¬%��Q�1��s�å�]t�}�o����}I\  ��唺/�pm���������ș���?�����_3A�s�2<�4�<V5λ�/ � D���0�(+NL: ��z���� ����4\	i���V2
�ǜ�|��?���J�H��!��A�x��O�Sy��ϕ�f����5��R	���uNc�k����RþeW
�E����?т������RN�����Bä�.���-�@i��h�ij7�l�:��6�����@S��z���s�/�dN5{�&�M�0��ie�)�f!kV�m8���n������r�>���pL碆�=���%[�J8A�4����0"�BX
9�/$R��L�Dc	�*/mW��_*'���B?{�y��8.?���8����KNK[8�c��I?���eo6�EI� �|��@ͨ�lxr m�g�]�����a�a�s�lH�9�#HL�<;~�_Z\�{!�s�� �K�,�I��Ϲ�[��3Ӳ`�Ͱ�Z�e���s����d7�d�������{F�1ɦ��Щ5��Q����̿c��y��:Zp�ߪ��¤ɓ.Zpׂ;��q�)Ù��w�6�ؖL~�R�'fN"~])ˠK8 �q��a��ٿ�]�͇fO,���k�+������Y�0�!��6��5Sq[��@c6*��}b�)o}Ѹ�t�d#͔%k6�I(z	S3(KW.%�xL��^��6Q�VsQ4�ׂ89��3ʩ�.kkH�rBݜ{�xUt �͒�*<D���^[� �  �Y�+%Rm|>���-j���c�Um0��/~�EȬ*%�t�Ȕ��B�t��̱���Z'�jWe����Y攥�.��Z�|��֪]�,�r��k?��1A\$�]���ح��+	�\М������`�_�F�;����4�JUOJ�(_t%�'D�g�M�2MC��؝"o�����^�|�K^iO�F��c�Μfl2�M�}5���˂�Xk3K�a��U[�&�q���������E1w��VN<���6�̉d;3RK(�Y��$U�H�X��E�%�l��Tid������u�����й���F�VQ�8�m��Tm�������Ǝ[�!��	�4zh �V�U��������)>����D?B��¬v/}}�=��A�;���>��7�!�W�����#6'��Bm|��9Pko[���y�@��+,�#1a�+f�k�� R��y�{�5#�a� $<��%�Y��VUJ5K8Lq�ٜ�(e�WT.F��?gn?��iܑ+�dS����շ�dRZ���C��8P�O���@��8��^xi�����Z�ro���ݚj��y��dr�jf6��a�Y�C9f8�����gt�J!㣥4!~�	0*�����͇%F�|`!+��uP��Ϡ�@��_*�a����p){[D�k���ԓ�V�֦t\ȅ�moڠ�|0a�٬C^�	E�0%b�V�l��O��F#ڇ2$��n����%�O�ܼ)A?����2����]ˌ�,��?^3�V�����h-۷v/%N?k��9�� ��w�]��{�}���N����K{{��{��e��Œͺ^��TֱA�J��

�]4��;�R�:������ɫH���l*źb�Tr�a�hݝ���S+���,6߲	y�񚄴%;d�UkBR[\��mE��/Eܨ���c�ir�J�/	_ֻ��6����K�υ\�����.W�'�L����3Q*#񀟌�Dr���t�R���|1T��C��Sh�oξ��B=K!���&\��;�Nf��R2�ZD� �q ��0����Yw�%��Y�J��+b/+����/9��O��yC��_�B�q�R\�똓�|ù?C��ZG��w(g���N��\�=�9��bn8�	H�S�_���޴��#��|*<���}�q:��	���K�6.�tZ�@&��g��U~�Qio�T�ɯ5������No�^{[�>9�F�Y,JM<!��V�={7�䒋�e`&�a����SO��5�����{�m#���J6_�g�yFc�-ӏ�/��6������A���~�3uH��+����d��@Y$�Ql�u;�SW�P<�j��#����	Eb��B�I��IM� ��aɤ�$^�L!+�X��c����A��6*�AK���� ��j�J �2g\Oڅ�U�AM�f\Tyd=�X�o%��B��k�s��À������Q�?k���,4r�܉'*��7fv/�`ʧ��	&��#)���.�0�����=k�Z3������_��SOy�~�!:T�m�j��e�/��!3f�R*ߘ*�_������haT�LGt�W5��9�Ǝ-��8]<h_�(U(d���<%�$�6l��-�ƍ3Zv���t�2e�n2f�x}0����I����9I�[����EL5)����~�#��6-�8Zs�j%V9x[V�t���|ø�J#�;^K �0��X��ĊiɈ�:����W��nA*v�[e��骍Ȕ�M���[`�tە�_^x�����'K�~�9Wˆ� �-��X�o�X�<C�A�`=0椯z6}]���A�@�ˢָo�Ws.�{�t���1״y��1׼�s-���<�߫��P�����|ǯ����|��=��x�;$��X,$˖.�GDk9%;�5󺶾Nv�<UN>�4�y�LIC�f���C��o������=�h�3w��$�mWW��!T��#�K.�PR�.)�R�ʫ�ŋ$�s�(�X�����1ǟ$3f�f	���A`a�7Z�O<���{D&P��/��7߬ܧ��i�Cs�����W��j�_߸^&�oP��D���D$+�LR��V��rӍ�	e�x��g�#;7�(�Z�,%����JqMV3�W�O�GKw|�d£�yY�k哟��$�W�����b� �8���"�|筽g4���Eq>�j�6&����9�~���ܿE�Yč�*�;��<{��A�ܱPp�c�0�F��Aik*���D%���+�ʋ/>/�������b�����%��%'�����Y�����mwܮרV�b���<`R��!�/�lJ^[�P�lX�$�74�:^�Ԥ!ʆ��;���TH����j�Z��#�<��$��D�G ` ��Oa��ú�DYT���+,΋���b,Յ�^{P��x^_șF��& #�M�0n�\����œ�	�%&]͵J��"�L�����K.OrRX�4ΓS���h�q��_��Co��~U A��B��;�����l^���~�����߮�0+��
~���`�E�Yh�i�vߦ)݈������ޤ������n�F	0�ǀ�w�o�Է��<��E�*{�֬�t���.��Ȕ����L�SR��e�ڕ�a�:Y�����N('�C[7wʆ��RW;V�zϹ2k������������s���P���&7\<"���̝��d��#�45�����U2��F$��_��^����%��U�WH6�rE�����eg���D��w��o;^{��`q4A� �l(6)�>�Na$:B뀈"��"��h�9�q0��Zp�ݶp9����1OY������Z�F5���)��/I�8zIB����N�����&���ߓ\�[�Ѹ�i<K�M�-�|t�௢�^yu��[��u�����L�Fƕ
�1? ߂{�|p�U-�
��=���QHe����{)�}�yM�X����	���P��Ox��vO&�8�w W��r�a@���57Ա�I��snj#A�|�+_ѐU�a��?�����ʻ�<��?�S���'7���>&���$Y�f���V�p.$�tNV,o�H�N6nL�1ǝ('��?���^��%��O�o���Gn'�*�O�B6'{�>[���5��꒮���}�rһ��b�G�4��Q@���I��KV�l�t."�W�ʁ�5�y��8���Э�;���A3@ۇ�4��6���
Vv�8},�e.���ð�B B���{���-�&�T�B�����w�!����$!�?��$V�h�E��n���}�����eΜy�ӌ�%O��W���ުm~7���.+�ՐK! ��=4C���R�4������]E�WP���]�#6e9	�4���O�X�A�'�0���<M�)ꏡ\[5�2aPm��ތ�7�f�0�i���s�Y��y���/jH)�$���sP�xAa��p�z�ed�����
��M��Ϗ�J��wW�0a�,]�DR=���LQ^Z�D��'JSS�4L�.W_�q�������X����-�����G,��vz�w�ے���+�
��n��U�R��>������C%����HGgR%,}f[6%��i��N��h��<T�z J����}�Ta�nB8By�L`u6��f�F��z�D�+Ui�V�Tw�F�u�Y��EW����� ��8d��xp��J��qh?G����-�~�
�jK�b!,�PN��E� �o�����wϝ'Sg�&Y/%~p���f�'�lU�i����[=k����W�������@ɞ�Qp��E +��h�*�O^�L�[��� ߄C�1V^v�rJ���E�ʩ���R�-�g��k�Q9����?�i�+ <�[Ț����<Z_�җ4ʏ}�g�}�҈�y���SO> ��L�0V�-_,�T���;�e��ՒN�ds[��������F�+������?����YC#��46~;ٞ�XE��Y3f�G���$�QiٸV�ӯ����p8%�ׯ��֍J1Dc5���)�[$����u�2}�n��O~R��L�u�]��ll&�Y͛7O31�������$n�\�b2��-�8�*��9v���{�:�D�X�����X% ���u���)�>+�ʲ(Gq�Z?�A1.���
�;Ϳ��N������Zy��g�ԝgI��;C��5���6�}���F�G��>������9 �hno����`�?XW<����)|+�5j����JM4Z���T�P��}��0�V( v���j�;������w�Y��'��	�TA�Pv��i4�F�S���6�oʔ)�-W�Z"���>��ݥa�hy}�2I�;u.�+J1&���H�^��9�������_�DM��(��?�ח/���✹s��L��/�W���ҢL���|���H<�h8/�T>ho)�es[����ꦉ��=���5�d��Y��SNx�)2w�\��l����'[l$�8�I���eQ���� �-����Dk��PIh$�;��R!�l�тF�M�O}J��7�������DC���v���$�����rىb���-7h=�p�^N��?���:�������k���Y���n!����X5�j�3�ʱh�PD���|�V5�&��	�ٳg��F4~˲-�N�Ž�ڻ��HM�����)(6vߧ�y�{&��V���*�p� >N_,gzPn��n�����3��g?��ww��SO�Fv�e�����U����Q'.AX�.	�H��69���e�Y�HM]��Q�z�J���y2�gräK�ϟ[���__ح����E]S'����-��!5�<���2vLTZ77K&ө��<�I��d�Ƥ�i�,m���+�Y4���n����o����6.)�d�ZV�ղ)����%nX�E�P�j�x��<����(��s^Uƅ	K�x�.��LP��f��a)�sr�)'No���OL�@$=��&�)��o�;o�A����i�g���H�8�Ԟr��^j����4���L��1�޴ȵ�u���/�Ɂ8�yA#P�� �4?+�փ k�5J^
�4� �|fl����~&�����m�������Z�q�o̲���e��ђ�X4��_���g��ǔ��N��%��l�[6�4���O�|(!�6u���kecK����d��p$"x�O�8��t4A�����_����k�q�G�|@ҩN	�Ҳb�bY۴LB����0ц��	��²is�L�eO9������Z�������i�?� ���E��ԤZ6<����M��$y�:O�R_W���7F��DB�r���fiK[�R�Ԍ��lA�����P$�)鍧�K��;S�uǥ�3R���-���;�'�ߩ3f�_2�i��6C�M��<���8uU�7���c�'���"�L���:媫�ڂK�@8�s�_t�E�\�SM3C�T�4p��N@���~�ܔTF�	�ZQ�G��xs����(<p?|�����%|Yة��T�d��l�{����\z?� 7���ɼZ$�|�C���l��j> ��;���
�Y��"�Բ^
���ջ�n�V
��,[�$;M�.�x�I"r�P�k�dR����'Mn�l�]~2�4�j_�,��y���������)�\V�z���<)���	B"�e�<i���]�!���S�5�
����o~�	o���_ %z��g��X���e�Z�5�bc���J��U�I	'�?�X����
�!g*����"!���:[�q%a��J�q�����~����K/���~�kFr����3.��?�W-�j�<��s���*9LK*����os(k�ݾz����o��,[[*��GT��M�lx�>?4dӢx>P`���_�܁�P�cn�u�*`�Z������`%� 0��iԈj>`e̕�c@��8��s�OV =�q^�!�,ɑ��mfB��"֞�� 2V+��t�2hå}l̾���p/���P����?�Q8�n?߳,`��L��1}����Xs+�.�t�GǬ�%^#uu�d�]��#ߪt���O���n��]�j�W���{�����2|��O�E�`�Q�	چ����>��j�(6���n�g8>���+��( �w���i�(����v�M���ok� �C�fX3�j�OooY�h{i��U1/�HDk�G�Š-ڹ�x)��AP����+�B�h��$H�
V��z��,ި�%���K�mG�Ux@��Mڹ�y��k��Dr�r�-�ӌ騂��2}癚<d���9T����0�PL��'>��>	hWW	.��-
�����@��>p�* �mp��    IDATk��&���7��u��h��#���/V��^Z�p����~��G�g����̾"J��s<[ȭ�B�%�k���?�#t�$S.^�Z)+8̧�|�߄)
������gF�|?sl�c|�#�Ep��1��fT	&��a��B�{3G=Y��~�3�j�ܴ����~�z�Eۣ��+��$��3�h����c,^k�d�Z��駟��k��4���� ���4 "X�x��u��jR��BAM�bT˰����G��Z$�m��R@A-�E������\Ahd?�O���_*Gu�V��������z���yN��M��p�$�����&��j/_�g-SX�4,M�"������ |��!��ZrbEdQo��Z�L������7ARm��ל��@?�1��/|A��=L('����� <��K��I�:Q#,��s��!b���D����b>+��wh�}�@����\rnY�����!���uڃD�g�P���<�W���=�����X�p�V���������ϗL^�\��ˊ�tP��zݖk��|Nj�Q-���~�.�K#-�)��`�B8T�����2��U�����S��4���4�7;�w�v��ш�� ��'N{SK�
�lp� �� �X��}H�k�������v��m|f��� �;��wܡֵ�a�<����r�[,,�
͟(����O5�`��Y����f��v��V<�=> � ZWR�Ǭ�� ��������:JKD�]�|�w��P�
�C��a���Ϳ�#���1�����2��Ĳ�X��e�Y�"�3�m��u�^ܯ�c��]q��p���,�j�8�~40�3�@,�El�j������6ܾ�����I����4&?Wt�xE��=�?�գ��}�A���ϣb�?��(�(�or����F�F�� ��@��}~�NZ4UA��������?c6�Ф��*Y�80�o�k�kXn��?B��g�ؗP��?`Z�6��傈�s�'؀�H����&�/��BIq�Z|�%`]�u�����1c�j���B�h>~���a�U:ۻ��������t�Ι;����k'��Y�.6̀��$eaqF�w��O:7���/	���-|�-��P�;X��@�-���>�C�@؄
p�QI�H�����.4w^�܄�����4�j௙����>�8G�>�������i4Ž��{�/�9|����g�h������_\��v��m|�4���t�w*M⃿s�;%��
6͟=�%C�ǣ�C���?�����/ �|&��M���m("�Ц��1v�V� ʤzJIZji�M���ʭ����b)�7�2*��N^#4ο��d{�r���s�ol��i&��AZ9�ɷ0N��i<��o��,�dq�!��ބ["�z���y���8���P�װ[l��4���?�q�h���p�M���������5ZY�h����\+� J�2��?������Qee�.��(h�O�~}Я�����?��1m�/���"�������1`6��2>ބ�Y�������-�������7�Z^6V�5�r�+ױ����ƹ�?jK&/��&�m���<��o��k����w{�v<��Y��%qY�-t~�>�[A��Q��ĩ�B�9�q�.^���M�/Pp_U���}x�,h��q����ڧ+:]��1�o���i�����RS|MD���$�ֈk�u���LR"���3Գ��7�Ǣ}��њɏA��e��r��ڱQ2P��	U���t�6����iS�6�xߺ�Y�$���ri�����m���9�y�ʼ���{�
V�k��_a�̝ss2�~i%�f�BA�0p�T�຦hT���^��_mCb�
̴R]_/y"��!J��x��L��X\2��d�"�0�D�.@�8�[A������ΔS�}���E�@���h��>��{6.n��z��WK(H�y#���'Ml����`��U+��'#�N��f���LHl���3��k��i5�xȤ����󀳼����m�vaw�]��A��A��A4R���&Acbc��I�Q�`��&%	b����ԥ���l�;;����{��s睻s�.;�J��������k�-�9�9Ϳ����!%�kF}�9>�|QHϿj޼�_�I�%����Fm��%�5á�N�ܔ�ɿ}S�?��6fa)Z@בE�@�,I(Q��H��Gs:�cZO�h�,喖���%ʫP*Z�R5�������Th6]��+������V�v�ε���\�/9|�}F@�n���M�(�v��~}Y�M4�a��Z��V��h� �Ƭ�F��|�
���袋<�h;!��C��j+�o&|xV�}h���F�����^� ��x�o4WR:]	{�4ք�s���;�����O@��Xf7��ȹ���6u�5����%�R�m&uX�Z�l.8�� ��p���eZ[lm�z��h�j��?_1�?�2�P�bs:ϱ����8|Pr��ܣ}����O�������<շ��� �������LE7L�?�>ǏF���u���B��{z�����%�ܾLʎ7��	%��Q\X����FC���9��������8�I��;z�	�����J>�s�x��~��i#��8�CŞ���yS�X���T�/4�UOq�\R��l%��$y�����Z�>K�zp	���A��������ߠue|�AAP��R�j�~S'�%��t�3\�
ȎMm�;֚���v `b��5Η�#�#��N4��*�������3.J��b�wliku�u��Ͽ���xĴ�"���hA�s9�3Np���|���M����#m&6�M@<�����,�ac�h�x�����-����I�!L5�#��*��[X5���+Y�J�}�m�����3�i�Bۉ3�8��r�EV��]�_p���C=�?�Xdn���_�MH�(�E��P�f/�'M>�jDT�X׏�n�{������Xo�C����
��cy�0�^�Sۭ�lh���'2��9��4��E���/�����V�o0��t��5{����ҠK�ġV��q���P~G��b�+�k<�(MχD9Gswm-�,^"�Z��ʹ�{6��įJ!�����]��L.���J�5��H�/UҞLv�)'�e�����3�-�"�'����"�������6���o�Ǎ�}���B�KȺ���M]��KqX*����v��I�Xv�B�u�l:���0�XWZ�)�c/�J���8��ⱎq=�SO�	W�Y6h����x���� "���O�6X�B�|5m���D9(�wSP3��뵃^�*;������L	��=ے��׮��]���߽���x�0k�h�T�|�	�ٕW\��>p�.<��q|yv#Գ��R��/�'��M/���2��V|~�p�1�"�?�"cZAʋK�/�����h�$�G�c�����5ݍ�JH`�C2}ϦS��M}�?�y����4��1���=��Ϝ5���o�����O���Ku��\RB�0;@����o�Cʈ���`1�/n4|
�Qȉ�Ʉ�@M@f<�F�?ׄ�)��v��ϲ9�����Vs�fq�fF���Yw�z�����z��{�����Y{�X�O�y��!;��W�UW_bϳِ!\-ZKe����J��s���iU���W�3�c���t.�B�� @A󧄂�q�#s�5������(�&;X��W_I֬(�p�\@�84�,��]2ӳ#l�7�c#�����*����>��@��G-�O�'l�$�������R0�s-�P	<�/`
�#h�0�ͪzVK3g�x���fq��c[[��f"r�
���a�v�y��C\���t�Ig�t3�����͛�l��LUi4 ��>�!|�{��@�j(e]��ߴ������F��JR<�1{�l���7y�>ז���j���3\qՕV*��b�h��p��d�z����r�Q���5=`�r��U�[� �f���v�yo+��V�T����A��0���Wӓm�u��KLOp�ui���5�`�j ��8�\o������̈�\2�4V��I<�l�/�3~��j��b ����<C��#A*��`�
��8��C<�u��h�D�� �)W��#���O<a+W-�r�j-�4�
ax)��G�q�-�jub����}���/*;Sj����zՁ6iR{�$
�ļ�y��/U���@���뮻|�dV�V5o�6<1�h&D� �|��ޡ�?	;���aƳ�Y���Ѵ��n�lB���>��������L��'���כZ ��
Dۭ\��L��J]I3�U�͛>����L�ٝ�ێ����?�a��L���nV�NVP�����~�%�U�g���0vZ߱,v�}�9}6ָ`�r�r���Z����EK�BG&�;{��9^�eŚ��R�8��c^k��q��M�p�Jh���6))8���k�y������B�`��ϴf�ђ,�$`+�'+fvg���=�kE�Դ�JH��q���/����5�b�`}��}r����͜i�����=�2hȿ��/] h�0�u@���c�Q����3�\��뼪'�%,b����Q����k"ph�'�P59�c-��P��Ѿ!�����nSuJ�ͪ�3+�Ղ��^Ye�b�}�Ϲ� M_�ﶓ+#�[�ol	lP�2#�9�����VjٶֿVB�
�$����,�3A."-?��a/J�b��aQd��5>�	篨(�Y�V6�����7	%�1�|	�gǲ+�{Q���9ԭ 1��׼�Zr���������f*c����,C:CK؜�E��O��Z�iߘ����Z�К�9�v~��;}#��}@�6�LV����㏵r�`��m����k��8y�n!���v�񯱝v��
�Р�ʄt��s]��G��u�8���?{�w1��5���as���FĢa'�X8��gu���6�O��]v�e��?Z�g�j�b�r�\��]�Q^e����͟�J���?{ι��n������V��ץIR�: ����.Vi��c.m�1�����V�t!.�\�k]+XB R�&i��˾�}�q(n������jo� ;�}O�q�o\L�Y4�>�o|�y�˦-C~M~�=�Я�_�<�T��ε�Ge��q��N/R���ݾs˷���V�X�q����z��74�R1^��:�����k��bi�2���X��~�z���V����S��p¤�מj��� ������pg0��'�OO,�R�Y 4p�q�<���G�g��g<�����(�+L	�s��$��IH��ў��
GWlֶ�ؿ|���:"O�5W�\����W��o�w�� �v;g��t�s�5���9�T{F�y�����
�l\�5���㙻?�s�*�k��M�Ԍ^ �Ϛ�?���8� @q,���ԱT����:�q��g����}�����}�q�{��l�vKW
�j�2{�
�5����!�r��'Y��SՌ���cg���aͲe��%	���	�1s�w�z�����O>ڧ�����ο��gҡ�+���;���-�.��yOY_��\�Ժ׮��g@�kw�Zg��e,d�]7��;�Y���ַ�A���B�w��S,, �9?��3������cNqS.�)KRB��#�,q�Ҷ8g��CSH�,�m�N����-�	!��R�Z�U�V{-W\g����߸���m�s:q������sd�R2�[Ç�s�HX͍��
�l���_A_������l ���j���O���O�aq7����D8Wt���P����3��~�;q�����?ֱ�p��ҬH��"�d*W���Ъ�O�V�(����~�"5g�;�Ӭ4�o�}kl�����m��.�e�����T���ݽ�v]���~v������6�c�}�;߱_����'�
�fw��9�����!��������v���K=�e*vם��1Gf}�����g\��j�[�.o,���ڲU�v��'�\��ˤ# ���ڦ�zϸ�hw�Ue�}��x�����{*�&֬�����X>��a�Z�)�-�O��uLF[Iy��ʖ�>˖�Y[e�Yq�}���Y���X���l����
�i���Ӹ�뱗�~�ӱ��Ib�{�i~R�:d>�V�}zZ��W>~2>���W��ǳ�F��Haoq��gu���-$���4z
�3�{�����k�j����7�[�����i`�_|ћ��4�a���3�K�=kJ%,xƏ�㾮��2��㿴�P�͜��=;�i[���{�
u��E�ʴ٪�n;�����ϲt��~��Cv�w��@o���hkuBk��tv�SOO�Ɔ�5��*��]��k�=����k��w�f�q���Ru�E�\_\���A[�d��*��pq����������Gc����8X,��;��}�+�WZ8���ŋ�O�bO��9�6u��<E+(tT��4�X+��Q�f �3,��ђ���Gl��휳��JѲ�!K�z����T�Ǿv���S� ��Yi��W�~ɴO<P�ų�ʈiJM������g��d�>���[���O�����'��-�y�3oФ
z�#��z�OIg8t-��3Xԛ#�^�Bk��b��
�_vɥ����}v����4�~��&��k�-�6Qqt\�b�=���۾��bS�L�矟�ډS�ٜ��y�b-ֽv�v�y��򫭭}�[7}�f[�d�V�o�@fϙ���|��������o�\{��Re[�����e��z��}�յ��z{���U����]��?X�EK��+�;������c�|����BF+�ē�'��{�mT6��O⋇��vl4��Q��{���U��P>�=e�4����Wmr[���!K��<�kš>+�)��\K��������v�G$6BbD�n ��,0��|b�Xf�+�v���RSt��h�/��'��3k��o}�7>G�˗��%�?~�����X�ƲҮ��Z;��|�1o����󛥜�����I��}��uk�zT�BTIY�?��}��i�@��g���{�q{��w��G�	��>���Z���Y�X��O����|�������g���]0|��_��_������HMh���9��?��������Nv�uW��t������)'g�L��?����>�����l��%V�v{qI���+݁��ô}���_Kؒ�/���ooG}��s�9�Ezǝ�s�@5��&����n���8&�%�9kC��p�'�(sV��j��բѰڥJx[&kE���]3�y�b��h����I9d#Rd8HkDZ�f7}9O���F&I:��Yk�e�6z4��6�XJ��v�o�.�x�Y�H��͟��3�я~�Aozӛ�W�j�*��>�яz����>����m��=��o큟�eG~�M���-\�B�0��
Q:�b�>���E��)�G>�	�2y�����׾�5���s#譭����sf$����F�O 6k�v����`�-4#)��}ێz��V�5kWY��5.$hX�b�J�^���dE�q䱮ɠ�,\��#~Xtj�ƽ�T� |��g?���{｡v~�����?��c��@�r�nC���%� �8�˰��L��28d9��V��{���� ��A���}�a���w �7��J���d}lrix<�k`ԉ���l#P�(X�P5dU�Ҋ�c�?~z���������� �F�O�s�y��Y�{���_��g��P�(r�]v�;�|?�����O�����U���w��{�lmm-�l����'!�<b�Z���t��s�}�ʫ��z����^�%'�JK��Ϛ1���n��k���'��L�omi���n����暫l�=w7��#�����Qجh]���W�T,�C<��s�z]��YW���~�����;�?��O4��tLS�s��n���������8�R�c�m�m�Qj����Kg���њ��gCW,GR�ӡcX1]���,%�	�䟁2���ޗ0H�x���@'p�c��lL��
(    IDAT�?�K��(IP58}��f���۴i��+�� �i�8^g��e
�D��p�^~�e��>��5�>�����C=�� �����<��`�|������ͯ���cOe=�z��d�
�Z���/��?�Ֆ˶;�t��_�tv��CMY*�<s֌+o����N@����ϤP��M�o��k��%m��?c^��&Y�R�����1�%˺l�=��#�<�@L0Q"�/���F �����O��a2zz�{�v���/Lڗ��I�Q^>!d�V�+��P�V
OQ�7�T&e�T�J��-�.g=s��?)�7raK�'{m�[�v/�:�B]% ������Fxr��(�F��;��ֈ�C�� �G�����-���W�"<�M������W�}~G��-Ͼ�� ����:�i����V�E�����˭l%k�d������)7c��csm�=��O>Ͳ�V��l��η=wH�ӈ�JJ:_uǭ�~e��ء�$y)
I~������ra�Vu-��}�y���?�×�a3��̘1�Nx͉����y�;��mh�Lc���=���k5u�5�M����s��Ga�,.%em�8�-��]8UCMO���:�4 w�d���0%����2�!]	UC�-���U��� Ц`3�x%��Y�>�^����7�w���h�?�n�Z9
�e������{�5׸U���8�������> w�ֶӦ{�t
5����ş�/��gS�~A��;ﴃeR%[��E����l� �@w���[�~�Pr%e���n��ez�m��Lo+:w�\��׿�B�YT�����O�{��n��KG��BU�C>8Ak�Y{G�
�6�3������h��Z<�v�a'g�;&Mqg��������}4�~����JO� m�����;(����3�BMSZ�c�+N�x�>���f�j�rմe�L�R�lE��+�%}z��L�J�@-\tʇۖ�!Z��X����q|�?�S��ڐ��8|�͛WK��8�4���]w��0_(\�3ڇ{�\[;����+.�k�X���G�M��߃F����[
����>$�N�h�\.c˖,�����}�����w�o�Wڱ�g��S���6~�B͠�R3Z�B�����n��扨�&��~g#�'��5�J��\��:�.��"kk%��6���`)0�CC�E��~�Y������MQ�C3!i���������'�͉G�$i�\��@ �s����e�� ;��sN��g��-!]8`d��cx<�f�kc��|��˄0OYX�ކ-��Sx<�����7Y+q�'mN�$И�Q��Q��X��v��w�Ã)ثh�(a8|k�S�u�a�0c�������l�#��Ѓ���q��5�чɞ'a��5�F��cO>�d;�3\9t�X.c==y���m7é�.ϱ��ߙ|#��p�w�(����5���sN����w4mve��7���W��N?�4�o�}|�x�\��0���g?�(����9*�8d�}�;���w�B�D� B��n�{đ�+��	5�N��6!B"u���8�{�>��zp��h�bn��]�A�(�{0�C�q�x���E��C5��y��������|�=
�9߬m�c�B4U(�~��b�ࠏ?�S�[�M���:1YS�t�]p��3N����˗���w�=����/ae��^�����l~�����ӿ̐�s@d@�f�{5ΤP$Q=$xQ�
�5a�� PQ�
�i���%��jqL��S�AN�Ϣ��f���f%��d&�Ae��H	#������R3��I�fB��_��q���7�x�GQ'\?���ˎ;�8��ǧ>�)�&eQ(���I���j�����{͝�WX7�^������K��i��B6��c�?�9��W�P"XZ&?E�H�H�h�7��?�X|�T��k�w�fD��b%�ȐEA��T%�ap���KfS'O���V(B���ڵ���z8w|�����w�?�������0gP:�~�pSwE��3X��@�?ɠ;�s�?ȸ`Q<�����\����, dBs��s:�Н�_Ӑ�I��2�Z�L�6�IP�1���D�9L��E��R������{,�!�����D;xꩧ�+$���U�g3��lsn�|ˎ�4j6�ֈX'�
bwGwRwF�z�IO-�=��r��H�DY:^חe����P�?�u��x�Մ/��!*����N���1|�����M|(� �Bӥ\k�gl�L/��a��R���P��U6�����w� ���W���܅	<K=hk�@�ȳ�?��FB: c�τ��sf���K�O����1���dVk3q\\S�8h8C�I��\ t&�s9����`
@����4:i�ٜ[�ݲ#�<K��Se�e����ޱ&)������� i��ט=�u�{�4O�?���xF���El��'�7 �Eϥ����R);�f�I
�Rb�^�ʞ� 䂕��A\K�B��<#�f��c��N^P?�>��k�P8��b:NV"��t����*�^o�qo	�۪���zgwv�G�'U#�_�Y�˱V���:���L���f�5_���ٛ��f�����X0�zg�y�Kw"pTq�"�bw<�s�[vb͌y��-��ZІw帎��i�zz��@����k��aL�H`p=S���@?J�ñ��艐 H<�8�`�q�(:=��%z�����e�och���I��TEb�h���/A���~'YiB̕�Z��,v�B�� ᭆJ� ����@�q�-��c�T����9�������|��F��+��A����8�J����-���\p����U��9oٲeN� �!�.Ƶ)���q�18�ڪ��,�X��Ġ\oQp��W�Xv-7)A�/kU��h��2؎k����^8S�����?9��e�d, ���N2Syf(�M3�SVl���%tmů����E#�ߟY���3�z�į"!.a,� ?��\����%@�@�1�<�����K44�+bc��j�R�5c�U4�s�����+�����$ˤ�yZ��Fc��i9G|?�7�o 2��<��^d�����Ƶ����t�s���L��?~js�4O=
�+������
����c7��c�����$\{C͸�Wq@��_�[5�O@[��="K�-�t.�P
NU*߃�	n���H�}�e�fp'�[a(���A�j�["��'��MLw���O�_�g�/xA��V�ϱ~�Jh�M�=�;��'�{�ܱf�9k�շ�r�M������9��Λ{��7�Xï�~bs-6W� P���4����z�������2�!��Ŝ�Kۖ[��C��@JA#��M�	L�f���a�|�$J� 䑲�7�.��2�Kg(^�=���@��R&��c�C��P*�|3k�3�y."Ɉ�"�&�l�X)�G�Z����˂�r�eE�;�b���.1:�g2D�T��	�-������U�����������a�$�Q&�%uJ��p�4w)�RP
�R*bZQX bc�Z�VgΚqՄ��sf%�﹬����I�b�I+��%�%�X�/�q}���LҖ:FZ�6�ứ��� ��5�`��e�b�S$[j�{]�Q��1H�;�����k�}��k�����o�|�����p�KQ2^ԣ�40׺�K줓Nr ���?�$3�9AԒ�o��,$� ��K/�ԭ	���.S$���p}�x�l��WG_�E��T YB�d.��2XE��Z=z�(DT�0#�.Z����fB^����ɐ�V�G�Y��=�St�ش�x׎Ώ�0�;j%D86���SF7	�f�w+������6��ɒi%@�F�F҄���8@ I��uo��ב	-gd�o��&�Hi2����^��I0ΓbPԥb�/��͌��o��o\;�j+N~4�v��������!�4.�2 ���_���[n���Ϗ���	'��?�>��>H� u���E� ���p�O�k�B%YƙZ7�?k�+�&�LLKĜ����α�pl�O{q?��P�)����$�>]�L���P��l]W�RI�j���V"O �V[���L����������>�q.�D�
ԳC� ��19��=�QH���o�1標���My�c�&K��)��n�$��H���Ц_AIk,8q�rR�f)��j�~��Ό�ų�ŕ�"��b�������B���ȣ���[G�Gk�}>'A�"f�iA�@Fc���/�Ў?�x��hŃ@��T傡���}��j�r@�0�\�gĪ �\�k�h掁�@�� �i��Z�B�2�����
1�N}��A��k�b�\R�����O�aKD*�%$ejs9B�O[K��9�J�leچf�ҫ�}(�b8�w��>7e=�t����E!庶�:�M��Jоe�H�7��'��ߌ�g�\�M)�C1�|�{r�2��M6�&De���MY4�����G3�5Y:��M��^Z���2XEn�`���_�4�XS��>����$���_�����������?� ^P6��������~F��: ��H�BB|�_p����x�8�K"!��x!<�}xA3Q�W~$i�γG�/��WrO��O �Bk�H 8��K�-Yh��͍Rj43��y����'0K!n�+�)�y��J�`�,��RVJ����)���Vk�%m���-�
���rnsC�s���hj�Y�(D��f�'�\&`a��Λ�=��7���1��] /
��/N��z �OR\[�!phf�5���~΂���#-8������^,t M\&�g�ӟ�4l����e�������C�w�ԃ�'�ZOh�O>������
��K�U���hd�}������՟�ٟ�` �n?�n�kB��~���=a�5�r��w������G<;U.���K�q�G��1���=��8���m��b���L�c!�fU�y��UI�80���2N	��%�[�q��L%k-�i+W
V�!KUKVv�?g�
I ��M��$�������]{�uȍDM)@@J�h�P�"D
���w�ڷ͒�"���?g�PO9[Ўpx[�qlB"7(� x��is0DV��c#��2ɘ�\�SE��h��=�G�}��~#���黥5YL�hƸP헱!����g,�k�Y���a��)����:��g� ܧ�z��J�_�0������q,V�b_�tVׄʁRB�#נ�V�@2�9�nR�@<� E�i��\-���W���شO=�C�S>p�Y|���U�k�Vm��w�=����V�B�bm�f��Y;%*I�*K�:�g��a�w(/���=g]��XO����2��;d�y�1+.�D  8?q��2va��M�3�q�C���O�	�GYh���~�8�B���0���L��Ϙ9�	�̥Y��(&II4H_6ٹ�ז� Px�����pP��<��.���¡x�E�L#8�-�x˄	�F���_^�/�;�28cΟ���
\��g�6�r�\1��5'�Ua3�����%*ǠBݯT� ��b�E5ȹ����|�r*� �i���7���Z�f�U���Z��O;��8�Dˤ����Ҷ�������3@\�;��mP'h�:q�А�,S����u����ڊ]�կ�j]+��Zmw�'§�D�T�X����Ж����c�r	氖���'�x�+�̹B`����Q؍a(��1}�hMh�oV�G`��
��s�:�N8�P��2���n�ZK���|�,��utLu��{���2��Ln3�̖>���駟��R, w��WOc�_�U�P��Sc/�L �����e,�{�t��
�Sē@_}�.�Q\��=�� 8K��zNC&�8BD��d�i�şK�������_�Z�c[��5�nf2U˦�V.��i'c�{�IV*�[*M�i�Ǟ���@��5�O��Rٜ�R-6T*�50�+�T�h�){��Y��+�h����k��?��m�]��J�^�)�9��4�VHyd�Lr<�p�y	N�W��?����;��k�S�T�U�,m�&4�7��$��*!��s;��o��P�![�b�����قE�\.��D�;��C�SN���lk�v�B��tcΎM$�_�_ٿ΅��A��sbPP�q3���P>g�vz��{�s���|�Z�W��}B��?�K
@����]*�������6�4j�6'?���:�F/͚��lTzAsͺ��(�4u�g���/����@kF��^ti���(�_�g$� A"Kgx�|=#�'h��n �{���٩'m�j?�>���l�v���<CJ�t��Z�m��1�Z�H-�ݷ��Y�n��"�m��Gm�o��RC�*g���h���w,ߛ���Z��=���J���-Mt���[�i�C��d���Bi��j�+�B����ʷ_a���a��y��.��ϡ�at����;V`�����#�w�Cה�P��'4�7��_�(��g߽�?��&Mn��U�����Gg��5�kQ1LJ�[�v��Î��:�'��&�0>%6q<�t��ALv'-��@m&mQ��EM!d����أ'�V:p�4,�x����	��T��c	2�
���" �!�/@�˺�8]WB�ϤM*�?��ba�k5��e��Z��H8�&�6���&`��1#��!�3�ϡ�U���~�s�k�ԓ^m�r�����mmڶ;��`ي��M���e�mV,T����1c�M������P���gh͵Y��gK�κ�.�j��ҩ�u��ؗo����X�rV&��7��g���X�g<'�G�[Y� �A�-`]��>�(��u�㼟5c;kɘ�p|rr�Z���Ckٌm��L{͉����z�C_p��9Y��Yi�����|���F�>���ʦ�6{��v�i����=��k���^m^x�z{{<b�D��F*e�Ww���C6u���_��ӎ	��~DgP���#D���	Ĺ��o~�I8����I�
����ϕ���S+������|ST�P��w�ѵ��w��a`�������@1S8fY��.Y /�'*�*�����
J�=�/��"
(~6	.�d�����xw���NT��e3��}�k����J��*Ռ��v�Y;�DҥlҤ)�΄օ8|{{��\�����v�P �{lh�ZrE�Z1���4�c)k��]f7}�[��b�T�U2P��T! 4t��=6��Y/�5�
�V^���}���3J�J�s�8�^RV���.[��{�鹶�7�t�?T,��@�֮[o�춧�~���ʹm=��[o�x XF�O'y��}b�z6�͔I���iӷ��2���w�=��+v�R��-z��}\S��ށA�Z�e�r�-�׽�ӳ5�8���-��ވ� �����pCy�������/x���!�|,ir,����j�c���Oc.���{hl>i��$��<v�BH���c*�O�P�S�0�"�!v��z�N��K� �yLO�7�*�/��{Z���;#g�$�3���<�4E�o�R�>{����I�=���>�fZ�c�^��nX[K��������R��P���´��&O�/�io)YO�E��/5+�[&�f+��K7�a��a��"�ԁ��y�u�A	c\Q���%������2��>����m�f�>�kKY�e�[�x�w9�500d�m�mɒ����V�Yo�\v�t�V,V����[n���h���&4�7��K�1lםw������X�w3�?�y����c\SX�|�5Pu�?���/\l}�f�W��~�b�z׻  z���Hh�LL6� �٘�9��u�U�\킀�!�nEn����8uƂ���?6�v��f�c�޹��6�w�99J�Ҧ 8�x��f��`9�b�&���u�����t��9c���Ɗ�QB1m#��A4�^]�T+���X�H�q�;�3�v�%{%Zt-����
���N������'a�r�U���.Gٔmw���oZ��B�J���th(OC����X�0��{��Y����׻�o�d+���7�ak֕\�SF�	�    IDAT�����_�>ߓg`�E0�\�`�PY�ˏ�dt3�(x0X�KϷ_?��}�����Y��s�u�;x��l�=�س��vؚ�}�������v�k�+W��<�ŋzm��"�W���s���lOw��F���Z.�>{�e�|�u�Mm�������c�y�ў��l�"����	�d�֓�%K�Y��j������~�����v !�����y����L����H<�y��>��x�v0�C�9��scC��[��r�4"J�F��{��>��̝�hb*@�W�t2_
	i�Ҩ9^��|��/��:�,��U��}E=��~=��Gk��R%(�N��_^1=U�p+%IЮ��Y �h�T�:�9�N<�(�z�Tm�=�:�Z�gY��/:��	`$w��������� ��YOOޓq�����Ֆ�-�j���{�k߸��v��b��MLmE�RԍVI<���d=u�Q��o��6/����C^y�^}�}��f�n%�Ս"8�����_�mGq�M�:ٞa��*EwDS�(��g/.Xj��$[ݵ�֬�O��=J�ZM���{���|<�-�a%`��o������c{���X.]�%K_�_��#;����R�ŋ�@G�˶8߿h���ڳ/���~�Wgd�����?\�h��ꪫ<��+�q~��pΟ"]J�  �(�J�l���q�V��ǠG4�Nr��$��o�� �l$H�o,�w�e����˚a��S�� ]O���|�)��m��@�?q�|VuZ��)�ɲ��� _����	�RB���[b!��#�w���W!�
��5�,U7�v��N�לp��J�VI����l��if���0�=X�sV����RgK�����2x����P/��
C�V�H\%m˖���[�ۖ-ﮁ����o�F�����b���_�c��O~��W�r8�x���|�#���z �������~�=;�l���J�h�\������-���Yת^�d��>�i++V)��ӟ��-\�|�*���X9���\�p�V1C�Y3���|��V)z&�7�q�w����UK�o}o����D^�p��*-�pi�~�1^G�����(�t��l6x`�Wac����Ss�=6��Hӓ8h۪�7����? ��;@2wp�l�_��מm)�Z!���UV��b����/�ιd��X����,rBD������B8��X��Q X[��v�\��ƽ�YOj��#Z��F����G���R��R�;o�T�,�1�Q��]��l������9�
C��ɶ۔�{Y*=9������\�t�ޝ���{�X9+���0���a�������
�P�ǭ��B��5��ׇ�|Ya����{��w�XSO	
������^W��f�c��"�W�Xh���ǎ�Î3l��'j��Ht˶�ܧ�Y�J��m��N�go�¦M�i]]��N^�腭��h
�L�J��I�f�d��Km��w��\������Ͼ{�`��]���4����x�R��Zo��%{Ӆou�`C0�ԭQ�8����cs:/�¹3��h��).��7��V�o��f�% H7��T�C=T�×FkYr�rGE�����
@0 ZD�!���zj�E`��gb>w�K�)�A�?k�{B'��  ��L���r"J@�kp�]w���p-��~yQ/�u�f+�(4{ u�_JX������W*���%����jf��b���#Z����ed)���@��U���r[�R��[*I����c�D�� 0N15w�Eفh�W嵳P ?����R���B́�&��ŖIlĽk�&������18:�l��նx�*��ڜ�7�QGo�t��>���緿S��}��U=u�J�&��3O�׿�4*���}���l�e���L*k�\���Zg+��m���|��j-����"�ŵN9���j��{�q��a�c�N��x��s����#(-Sa�lZJ{ �R!�����<�N�����bߍ��f��W	��:�ی ��Z9�ro9��q��g���# }��|�߬)�G�>פ�3k�sE��i+�D�EMd\�H��C�C�1]�G�����p�|�G+/�<>�R��M����J���H����B�E%�s ��f�3BI��uPM	�I"��$y�9GFio��G�n���<R�A@q����q�E�\��o�r+��.�[e�kW���-זAY�5k�=}�1y���^o]��-��oo~�%�݌�\J��w|�~����5Дc���������[�\�?�r������9�_����6�×����O�`���ˎv��o��ӦX�2d��=��Þ���i���l۩����w��;ʆ
%��@3d�C�F0��DBew٤�+N��墕�!���G����?����3��(hȊ�Q��;�K\U1���#iD1���hq��@������ơ m�K���h��%A=)	`�U�
�qM�����x�y���`�p" ��{�zR���� �zQ#	3W�+������'Y���ݳ5*��y�н�
hᐸ݆'
�L% �?k�U:C�^A�'1ܴ%� �u��ט�g}0�c,E�$OB�����c0�(x�;��x㍶��)�^�d�-x�9[�b���-ז�l*k�C�6y�6��:�;�H���N��jU��t�Ͷj�jǯ���`fwv~3ߓk�hB7����N���>�.��ki�X�z+�����'6�U�8x�A�ٱ��i礡�~;X�s���J�\B����4O{�����'_G�� [���S�WR�X�������U2��#�H��[���}x`�`�5��.?�/-PU,9� �@q,稜8�����Y[�8��(%\+Dk��*��{��f]J J���)��
urj��֨k�������Oi0�.Y�5���(Y����ܡ����h֠Jl]���U16�����7�D��+�(g�X� ���1���1c�Q
����lp`��Lj�+���w�e�}yW��:m��6u�t;���m�]����^f��q������En�F�?g��������S0C%�8��'���:�u6���z{�[kKp�6X6ko�_�Y_���P��~�;U�A�x*��BaC�,��niܿ�6�2/�H�M [��9�3�w�^�:Ná�V*��ŝ˪�󷦕FmE��7���}� �F�����UF'Bց�����u���@����7@3�:rfs�"~���q>���ǰ�P�$X}���.r�A.��i��qkP��AH{�ɰu�ţ����M\���o�;�� �[7RR�sr���Wj�FM�4X&��J�HI���t	�ׇ~�)�%@��B@��(��ߡ�O?�u64H�G�r-T~�vE��E��nc;ﴫ
���p�i�{��ahO�I[�H�k�WR�ab�>�;;���ɿ��.6}�v�h�y�v�i'������!U�g" 6�SO=�� ~O?O��)ڇ��?�����W�£X@d������
4I( 4:O|�V����<q��`ߏ��=+�s3�6���%�� ��ﰒ�S�$��|B �D�p/�s� 7���zA0�9��>` �1ψf	�@ @'r,4��s��\�Ǳ�[օ ]��m�X�xP2�څʀ�E&?	��9�j�2��ƥ��$�zR8w����	�>��B�}���������哀���� M���>hN!!,K�qf?3�8��8�o�� 3?*���>��{��z<(ԛ��z�ɧ���g;�8��|̳��|���}�1i�Sy��|�������Γpk�ʷ�C�'K18�B�謥� Tڴ�^g������Kd{xm�G����9�=�����#:�J�|1� <�lhLB6�/���������9�n��?�(ʹ*�K�s42�wM�R��ߥS��U`���%��a�3�̭Z�1�k����3� ���h�h�QQ�P�3����7�FP��$�?��5���M&J���V3��Ij��+!�)���q\g��c�<)����M��Ki��s�GO�I9�c9��4�kS�f��u��(��o��M4��$%�k��օ�O~��v�]w�~���+Y�{V����gM�A	P>�"�v�q{;��cm���9�-%�2tt��=��S^.~ͺ���*�vL	��dF7��gΚq���~S�q��s�t~�'��htͿ���R��b�r�!�'�=��͂$n�P�+�8������C(�����a���� �Kj7�=4�K.�������%{lb*�[aS�V�{�D�H&|�xw����"`�?��^�Xjr�h���������@փB|�+*��կU{L;q�k���N"����*�W�e���RX$|�'X<	�'�S��寪Y9��y�������0�k�W��^�`��0��2ou|-��F-�3�{l%�<f��|�U"�'^'�k2uk"~�v��; ��׾֕;4*��ЩJjd vS*>�
��P<4���|~�uw��|�$	��o�R[[(3aqo�Q�����C�XXmI|�����n�9fk�xQq��c�ɇ2@�3���dx>��N]s�5�9�}��j��7׊�!XDlLg@��������29�1�[m��ix��f�% d�|�S�rK�Yw�$?%�c��p��E}��qȋ�q�^��ω鎀�8�Ѓ!�������6�~|l
��>r�J��X��1��V��յ�@��f>��H�c�%��أ�:�kn!9�%P`В#�?���<QK�a��k�BeCoK�w�]F]\�}��KC�N���t������S�=����'���E�/�G�F��<jxѲs�׆j��˨�<��4�S �w欙WOH�������{.l���}#0LƆQ	A�	�b�VE|8Y�4�V$��=I��?�s/��v�2��Фah��Ѧ�
8��B;}���~����}�V�lGi����Р�0Nd�G[4��� x6At��8�3��˓���Q��J�s���$F��s��Xq�����߯��$�����f���b�������D��3vs.kF��a�0��^z|N�L�� �5Ф���y,(�^@>^�̔�4p�Ԭ�@Ŗ����)f��P�m���9�=��W���$5�j͉�1V@��/��-��ZK�
�|L��~�(���u�?�/��{Ml���%ߓSc�	>��l��R5�lD�Ol���i�M�?N36p~,���ȩ��� G�L{q����Eb
a���"�t4&(�[��-�������8xd�5Z�5z	E���B>c#�̜�<p�18�2!��)�'�G��<v��3L~��㇫e>��蚪���̋gB� (P�����<�� ��j��<E����B�9�lt*jJI�y��x&	]Yc���"�D=%eFV!�s�@"`�.���l�40��1|ox��Эk<�Ϲr�K�I�3ỏ,(~���o�A c��FBIyc��U�c|f��	���,�$�����w�ynRKsd���]M��9*-K� O�F��C{h�j�)Z��Y����{�:�+j���F}��^2�"P�[���E��O�<�|U"�K��><�B$�k��]V  �s���K��gNI(㧴a���9����"�T:��	8@�8��?I�=q�a"���z�B�)K��~�[���Nn��-�z%×h~P���Pn4�MDՉ�A`IS��r�+p��\�����O���Xh.CUP�:��Q*&�w5=���i7����+ƞ��	sc����x���6���k��fb�'0�"U��T��C�Ģ�糁y����)h]C�����1l�Z�i"h��67��Xm�,
QͿV#q��Y]�.�q/�+ A�:cD������.���g^T�pt�o6�cO/�7O�J�:J�����	o���d����Љ����Wq�����6�����B��f��y.��uyv :�s�.��_~i�Ϻ�'M�x�y��K�9�Mx�����j���P~g��x.��b�C�I�"��zI�F*ž��y����8]��>ße��Ev�-��s��4��p�&���ԯ����#+T4m}C�F����'�7���Fm��i�	���8�e����E68P�����j�-Pa�0@4%�H��8�
w��y�������/oX�Ζ�����$����d��Ҥ���pH����qrj��\[N]�<7��	ϕ0�W�) �f̵ J��$.Yrr��LkO݋��YJ�R�g	<���@�����}xO<;�������d�] �:Áy�A����ȓ�@�B�q.�o�w�8i�|/�Cd2š�Z�::s�G��"p��-�_*�C���}�(����3O�z\���W�%���4N
`.D5SNF 
5�^�~�
�1���wD��(�A����h�A&���K�!h�ld5��si�V��1��,l4=ř�@���V્΢��rP�D�/�7�m��N�F��ܺ�k��ъ����_��X����c��>�y�<�( �U�8D��&����̭曹��&�Gh�P9
��oU�Dx ᙹ'�����e��s:R*��15%+�u���R3���|b��L3�C��,7�A�<����^�7[�zUT	7D�[ �Q#Ifq�ŦM�nm�>��W��/��^*ݩ<��o��/�#���=}&z/����b!!�b�<c,0�	�f�~Bk�c��7�z]C)[� �5��Y��@�4|i��6��r�rY ǰ��81�R{��K� &��.�f�� ���t�fZ�,�!@	s>�	����|��4n�A�.m�EEc^x�>
I߇����?~�[J����o t�K������;2����X����,XB�S�>�g�����EY(�RJ �
�s�hA�N��O����`=���f���F�'` I�c>�`��#T�>=!�*�)8��Җ��l֬�m�?�Ψ����CJ0�D���t�8�'"�_B_�@���W�ޯ��	��[���sD���#��3g͸rb�z6)�6q��e-�ZN�@ҦT����X�\O{�簨��T�M���a6�;��@1�2'��M!}'͟��YX�i���኱�"EkH��Oir���U$��;]W�%�CTB�T�ȱ�N\�8%����Xm"}���T=�EK��E;4N\Ka|�uUs߿��Dhh��H�_Y�������xZ���3�|�s���y�=.��g ;B*	���yF5o��ǪDH�"+ �
���!�<3>�I���M��g��)�Ce�1��\b��GF,%O��޽��U��Ο}Ʋ�S4��a�n�������-_��È��?/�j*��p��֐�{	I	,�X�|m$ٕC���=*�r<�+�=���`�(	o��Em������v�Z@����`�y�v�I!:�J�k�V[Oo�ggs�����]� ����=Ĝ�&[�D�B� �-.���Х�iaJi��ڸ�X4A��:_Z����o�K�u=	�%=���_�a�kSmI�g\��3��c!!��g��������7��q����8t���ԙw��́"� w���#׵��3]	@�g�p��x�N��ܗ1�;�y\�.^�[�B3�;x>@��Pj���0� @�X��VD���
5��9�Ѓ�"o���5��D	8�6B�p������h���RY���5��/<��e8l�����<)r�'��%�N��qh��E�tl.�q���d<j�Ak��N���'�n,0�5�1K:�O��ϔ)!�pg`��AK;�������B�z�lhpО�;��1[�l�ku
��s&��?J��̣.���"b����\��h���c ��౳Y�4���-�A֎61 %kF1�S��H ļ��@�1�Z	��'�%�_�Z�w(������[C7�p|r�z��H 0l~QE\S@��XY<��=�9�q��:1�$�Psm>WY*�z    IDATG���{�
�^d������r�yzO�{��Eiq�rR���֐��|�;�i�|�V.�?��*[��n|����Y�~�lR�?~��n������~'���e݋��w�:s.g�[#IiW����X�d�c�M�����[���γ��	߇	��������������s;����_"G�4L-D��������4�a8��C��K�l)i�yY��i{q���/~�i��f�$�� 	��l^6*��hhp�t���'�$j��C�F��~i%��ka��9Oe$TZZT�֭�$�44rT�P��Q�]�s��X�m*�I�%�7��g���6�(�ሿ���2�f���ҸD�	����%�%,W�Y�þ��h ��<���`���@�7�Q�9�&s�0S�/�Pv|^�!���Hg:��k�tnSN;��3N���/a��J��(Mc�5nex�V!�Z���:��J�OL���)�-L�@N��E�*a�g�k�0�<� ��|��x�=QVX����9���;����K�ٝ��/W )c�أT��n���s;o�i��15&�EO���k�w���� �k�Hb^hlm�9+P�m���Z�}{��&d�����}�Cd��qt������I���
`�|�1�C(� uxӄ�Ȣ��8Wi��% `�'ϮD��;A�NDY+�4cA��&Y�L�"ekSIK��-�������L*8�Ѩ�bQ�A�4�ҋ���\BUVS���$ 4��?:���I�g�5M	%���<�E�i���!�_V�)O|���xM�9�N�_����GZqpȆ��e	�N}�j��p-�c�whiks�v�i~.�>p� g@��s�~���}$|e��j|�\%<�ȘB����y������,��T�M,L��BHպ��ح��ns�>�nO�k٪�7��:�t~�;�����ς����3N;�.����Q�`C�}�����?u3��6}�ǃ��Cl���I�C&�x	�㚢C(`�$#͗ʞPI4{x��_�E�ЬT$�x�����$-� �+��&���*G����Ǳ,T�?r�/�C�ݠ�dxg /��4�wBy):������f���{�]J���%i��1"��R
�$�%4e��/1� P�ঐI�ב��8�l�(M_օ�Be1�>��/IIF�3��
VF-���-?�,>�S����:V	d�{�Æ�/�u��3���.��?�iT��tu��=�(e��^Ƶ�oPl1奧YcJ�"�������z�2��;���D��ڿ�Jnd�xF��`~(��7_dS&wXGG��9���#�sK���
;�#m��l��P��>���ZWW�_��i2����3���|�Ս��X�l�]w�ٮ��Z�2u���d����<�+[�n��n���f���vԱ�ٌ�;��S���;�9~�T$��� �f�V �y������W�8�BZ��IҒ�*s\tE@�pB5�fA�*U�J2c��3�8�s��� @������Y���L[�c��Q�%pR2�l~� 'c��R�8�oi�G /�� ����ǪSct	'#�~��$��;q�S�=��+��se��)*��ay����D�`n%�@�DH3�Ж�Tm Y�(i��ro��i0���ޑ�QLX�N�̏��1�'��e%�]Y7D����;�_���w���e�"o�@�&��Y��).^�eoi�GQl��0��'ƛ�ZI�i)����m?s^=�Y��~���z����8�;�'�:�̳�^�T���h7��U_͒$'t�������{��6��-�gLJ����O�޽��=��\[�����`��q�-����U�l�̽���Z5	 �� ��(��g_�j�0�p�X �����E"ڠ�O(��Y��}Y4lp@P�,N4o>�"�cC
X ��h+���V	�(-�c�X��!�@)^�s���@ı,r��x>�%@����#��Cyj���A��{S�Ǽ6�(t# L?��H(�
!� 楱`��L���C��Q�r�ATcƘ2�*Ɔ�e�'�n�B���I�$�D�����q��K�zi�+	�f���X!��K�j���lHn+�J~����4��������ʅmʂc~�����Ip��!�G`̭, �7�Ǿ�={�����Z�E_�'�>�}A&Mj�� ���i��������v�gy�����q���zH�VͿ�̞3�������?�&ɤ�ɮ�Ϙ���������]w�e��l��EV(�ͧh�ۇU�cU[�v��=/��4��6��j�ڋ8r�E�_�$���~^r>k���=�� �?]����\� �hҮ�[� ���D�R!�A�@6 �6�|/��84��4{�� dXPb
��9;ƞ"� ^X�S[�����pGp�Mw�N^7��s�cm>�͙c�X ��+~zG�LƵDQ-�=��8�ZB�p��5�ye�r�1��!�$A]��;z�.���X��C�^� -
e��7�x��h��2#5b�t�Kb��\�ԓײ����y]�J�p]E�q���z��}]?��5�=뚦8L���/� ��Ų+�m����@����xɋVA�kZ�RM��E+��l��e���o����ו�{�C�6#�3ʺ�`���ȴ���OHh�]��?�{�*%�f*������t�1V.��E���\�i[���V�\g�b�.[gx�;rj������,�йP�3�I�������<�T�qj����7�KCf1�)�bt R� �~�3A4n�h@y@����;�	���U5ZK+���}i��>���3��{��#\�c�5[���ϳk�а��F�g\����b��������v���:4�l�XQ� �;Vt����M��jn��-?Ϡ"p��^ ��h�oE���s�K��N�g�o�%̽�L��M{�S+o �y_��~1t�
�y�.`d�# ���
�'%��[ ���Qx��|w,����σ:XÊ��3����}���`�ux��3ԟ�_��m�ݶ�i�;�g���"����\���y��*�zM���>��K.u*k��.o�l��Zص&����	M�t���\w>��F�?���g�W�{nx7K�.�g?���䓏�je�V�Zl�{�C͕T��u�ڲ�]68d�t���+��pL�����ᣄ���S� `Cv�a.���tg�Lhmti��4mD	iʘ� ��� 0c� ���f( �}�'��Nc��A��u�h��f)��}�B��0���1B0�q��b�Z�}b�I��-� ���(ʉ����k�D�W@�� ��;B� ߈�r�s)�|��=� c0�Z<'Y���.��� o���%�'�P�=��C���R�����o&b������{���w��?��2����p4�{��c�QV���>�яگ~����e�w� hտ�˿�� ��1��S��<�����;�C��Y�O�y����\���6�_�g�Y`����.��N�����������������hNa�U�o��Wv�y7{�{n�L�b^|�~�����c�R�׺V/����\��n]�-_F��6{a�:;�����x�ob6%�ڕYy�%�x/� �x�|h����O~�V��E�H!~ ���E�p=��j�9*��DE�<p��@y��@Bh�@(��P:�g@sAh���Z�|T����#@u�<��=��=TE��Z���O�TV�h8����|g��;D��S���`��F�W�NƇ�� Tm3QE�0WC>��������o�9繘/���،3�@x0�Xq�~�G�Y�ԍ����q/jN�Ys��P��=h��p4��p�ui��ǅ�t̖Y7�s��Ϙ����v�[|%���͚&G��o�����H��8����+���ڡ�c3fN�^���2�A2W�����-�r�Ŗ/�[�P��|쟼�iw�:���sYT�4��̪��c��/t���4�Jp2�������h��>km�ط�u�w�V.���e,�_k�����Z�Ζ.]iUk��K{m���eeX��,�h���7|SJ�C{@+���˜&��i�h�z���XXrk�� /�f� ^�L�C!�h���"U��o	�)�����������[|��Y[��u#�5��ⵡ"���~���M,���c��������\Cxa�J���-��y@H�G9n���x��k��V��Q���S�;j�uy�)kQ�g�y�x��!�'�h8͕H)&��-���	��	������ܷQ��%�K�"?��k���~�aW�k��C�A����(���J�͟�_��9{����C���۴�s���P��R��E֞|b�����_���d{׻�<��*��>�9[�d��q	>���c���ZҤI��w]o;n����`?���e��T���k=�~��,؋/,��]�mmw��?�-^	&$��~%K}�c��s�=�Ԣ��E�H��;��/[��ə�8�F_�`��I���|��L ���EI�i��t9ͅk�q	�Pf�d���Ikk-bHQ@�6����; �u��I�S<~[Z��{���=�??�S�9+UVL|��P����!h%��c(���z�}���a1��b���Z�2����\>S�#Ń��`�<��(0h���j�!�>t���H'	������׃�蟗r�M���;͹|=��1�>ڵ|.�h$���ކ��j I¥�3��V*�����ȦOk3��k�J�z�j �,�j�y�X_�Vuu��g̶SO=��i
eOo�֓���������[�\?^�tG~)C��?�Y�/�]�ٙg�n��>�z{�Zo�:[�f��^�Ԋ��X�
�P�����ޛ��]����Yg&$$B"�B�w"�Z��IP����ź�o�׶�����V\��KMX���(UPA@�%����6g2�Y��{?��̓Üs&���f�����[�����7R��n��$���]^���Z��c�5�h��[5�Ź�lX�9G�K(��}�r6i�*�`S�v�J<��^��xnv�h�C��܏�b�'�h��{	E#I��<�T��V��'����u	%�8�ǻ�X�����L� 
�8������	�J��w	͋�8H���w��%�]�KBw北�:�����d%j�c'&�AQ;ʚ�w�}4ǔ�@��Dsƻy"�~Z��0���N���(��yz���������/E-V�� ���Z��S�#ʕ��E֘�%]P	,ٺ�)۸i��ض�JղM��[-�����lp�j+�Zk[���eo}�͞}�U��~�;����l�#s�h�,��_���
��w4�} 6p�Cgۻ��v;䐩V���y���l��uT7������������C��N{�2����>�X�;�0��+�ʿ�Z��7����/���f��6��s�Øwf#+kT$�H��"�A��7����'ϣ�mi�Z�z�84��^�v���6)!$s_����eE+�~��������VA���&ca0�H��#�� ��3h���w���u�ݩԂ�c�'��X�`.8^�ɵu��+s�υ�������<��k=h����]�G�:��?~�;��W ��E3����������G��k\Q�����̄�rX6@�Y�YG�j+W-��+�yC�O2)UISV���u�y��c����`9���o�b�Q���V#�Ϝ>��ŋ_�8G��5�|��Px[3��dj1�ɋ^h/y�mBg���)[�z���w���k���-�-��ڬٳ�����{�M�p���¡B�P�MY}6�e����͆)Φ*��/�C�A�C+��6��ٷN�H�i%[`  ��x�7�V��.��K��I˽����J�����o��d���w���v�W�X�I8�z
���9�o��OE�$�~�Lڲ� e������" �oqss@�#�j�K�wZZ�Z?z�V��-�+Y\�x�Ю��s��Oi���9�_,9^����Z��U�,z�}4�d$���9w�(Ǘʡ�&3��L:G]����Ю&�p+�?������}Bg��c�s#��[��=��mdN����E]d^�r�V�^����,�e˖z1��g�9�y����̎:�y�7���w����Р�}=�}���;7_w�������P���f�/P�=U~�$���KmE���P�3��߱���cƌ�>�^�;���l����YX�~��}CSo?�'�E����rE��B=y>ORK���QYh�W���?���;�/?@��wh�X�y�X��CDE�rs��CWI��i��(��	�h�����|_�?�'n�g��Ϙ��V�Vi쌯Jr<mc%����s��BSS�Ɖ{ro���+��9
�9��^s�8�.�*	X渝e"�wAc幜���I�B�B*��y��Z	�X IK�����Z�\��|βD�O,������pP�J-��0�����)۷\Jh�&�ߘD��.<�T��h<��ݗ_� ؃zn�(� �v�*�%�O�l��vt۔��G`��#��b`����Z5�wt�����?�����B���'��?0�����.���)��w�PŇ�r����7�ѝb+4�����+&tǎmo��lHi�L:M+�� 
 ��[��V�U�`3�~������4�j���b�1�<<?��;�#ԏ���R���� Y���Ȋ xV��h�h� ���(�#\ �����w��g�TbB��8+�������e#K�f���bR�f=��k��}��)u\�1㠕ƈ�!��3��zH*zǆg-	LCƖ�b.9��C(sՐ��J��J� Z�"Ɓ
�D;�7��:4s��o~SO|��P���t�Ӻb�.������{�΂mZ��K��ё��M�b|�?�Z(��1ɦΘi���\���~���m��-�t�I�3����+h��+%G!��Zan�3{�t��"����c��;|/֟<�Q>x���e��X6�	�lGֺ:����R(��u&o�����?��;�Q<;:r������>c��nY��+��ߦ�c�[� kq�c�R����?����d�׿*&�����ʖ,y�^�%v��G|�]w��ݐؼ��ԅ��
��G�v�-A&�q��N���zQ�@�I ��ffa�0
��w�$#�k��.@Ģ&I�Qug ! _�HBR�H��
�8��1�t��3�q��V4Ҿ�}ėJ����:V�q�Xm���i�����T�&����g�4�'Y��	�)T�XT�[IZd�2~܏yc���/��a^G�S�Z;�Gt� n�e/{Y�i$��G�+k��^��C����%!�(%��sϱri��{�~�*���\&� �
��ZMp=��'b��Cմ�>�X�5k���6l�b_��{l�A覰,����#�u�%M���.�>s'kPY��Ε��P�s���<���ʎ:�9^I�=�N�c)�LV���ݕ�L6������ZP?��߮�;#m�IS�~�-�|���>@cp���*Ւ�\+S|q���I���|�	�I� 2|���x�� ��-FE ({Pe��w���� x��&͓{ΊL@!	Iڦ�F5o��`I ڪ������Pb�Ҍ��І%(��c�S<����Yisc��|��u��[���-򪬲H�)�ڌ��=O5c�Y+l|��f�'ƛ����an��5�B�C �@�ɪD�o���܊���=@���*�����P������������[b�u��V�Zi�6oXo}=֑!>�b�r�i4M;r����J[-3ѦϚm��j�j�
�}��k��ǟx�)��4���E	�� ֘񮪃$�]>1/���7�@F@��ɜ����#�������p-p�`��g�Ppq�[\�#O��m�f�*W��w�C�W(��UK���������B���>���F��
�;�x�5��    IDAT�B�g5YV_�R�/���2�/�i(����O�����^;Nk @$������rN㚊��Bi��(0�f/�Ţ�z"��De�*_E�x+��H�q�𾀓|	��POT�~W�6ׁ���2�5`�;C���{_���~�O�u%�>��@	2_rFs,Z�֔@a$��Ɗ��'|�o*�J��7��]&�c����r�s����]-�s��'�Q�xY	����?���=�[�@�M�r���w����趘���Q� �TyЬ<d�V���7[�Be��[��'/��CCUO�*��Us��9G۔��:�wz�_�p�=�d���!l2��.��b�Xrq`�LD�%�}�}�K_r˝r�u�]�E�"u�1��͘8U4y���o���PV^�*�?)��P�A�w�'���#��6�g���)�����=>��t�~ܙ��ģ+ X,�P��j�] ��OX��~��C��Omj 0a�Ӳ��f&���}��"o��3�i�5�U��X%�(�H}b�q�Qy5�V	e���`��,P����Uw82.� ϳbEȼ�;@�s�O}h?5$G� �|��/�k�\�Uc)*l_9|���i�K��&驿��#��
��8w4:�� p��\��^�U~�VI`Mh#�S���3�|�u&ڌ�#a�Ԏ�Q�'ϫPN �P2@|�ִ4����J�h�D��+���s���{,���Ƶ���c�ufҞ�J���~���8 תVM�l03��3�&M>���i�6��_���VZ'J]RZ=r�֚���|<ק?�i{��<�| ;�r.�k��}�<� d�3�Y
R�<d�X��4�D�|N�"~��}),�5�ã|�7B����Y	h���}*�g̼�L�j	��M��W/_$9,���31 VtO�P ���*�aP����������y�Q�i7oݭ�U��I!ڠ]��$L%TR �������� ����DkDp����y>��B&�@����;4Gq�,`��g��:��Q)��V�R܋��Se��K�_���g�]c��͏S#�q
%LT*�;|(�h�|���YT[�8�����P�*��5���fYc�J�MF�h�N\i���M��%��=�X��
�][%z�K�0N�Ԁm��rV�5�V��-����Ւ�,� ����TΪ�iv��ϵ��DK島e�v��k׻�c4�����?�'i1�j���O~�֬Zm���7����~ʂSߟ��1�Þ}}�k��D]ʊE�ↆBX1��I2����#���Jz�|�O�V�̘9��o���_k<�}����,*t.Q�'��	��K8�Ɨ�$c^�b�[ȥ�l�i��f��|i�, �8\����1�i���f�������s��sU�+�CX��N���1����E�v. �'@��@·
R�H��X�*7�3 ,q���� � (Y ��u�w���x
��DК��G ǽEY�V�C�Z�[\9U?U��Z(���������{	��h-1?qKF��|2��sJpKH�* �IDOi}J�ig9�{Qh��yN���i'�`��+C�~��c^�����ͤ�����A���?q�A���i�7m�k���=��S�'YJ�kY	�4Z͟{K@�;DΡ�S���N�(��0'�7��/��/�-Z�w�Y�A�Y򱐕BJ�N��)�(7R�5�T
ڧ���ߊ���-�I��a�g@��ed��ؑ�zh�f�6rp'�����l
�pπ�J5��]K�KE�p��.�f1�%\����z��,�&��k�+-��%
�N�)�x�[	1Q^zY>\[��! >��w�j�tہ��~��k��ߧ6.�)G�@V`�؈;����A|/ �z�
�JK���{�ΕI!�����R�RxX#G=S]�%]��.�x}����x.5�܃:Bg�q�k��r�i������W�N��.Tm�6�τ����߶�`_������K�ӹ �{��+�_�_
��]�� �1g�ׯH;|Z̟�nY�Z�4��A��9m���8vi���@5,�)Cs�j�[p�8O ��	bT �2����F@j�6��9)��'<���:�Mh	���L;�ԤM	|���:|/� ˃��9��:Ց��Ε�(^�Rڹ�M��Oi���j {����3~�����������v�Y����x��4F��"S~[e
�X��Kc+kP�1fXr
�%̹����@V�"��%4W$F����<�-��;�z� %��8�T�Ҁ��l��ֻs�u��CA=�\����;X��G?�&O9�JՊ;|���km��-MYD����h�I�/TJ{Y�1Zl5s��B�+|r��}:L�p�D��ĉ��aǡ�M`(��aއԑ��8���n�&�H�x�w��'�$uК[���~
��EݼM4yi�,8w6���ht6�6��G��1�h�I𝀸t]I,��2��'�]i�a�,:������������g�<���qכ���5��[�RG��(�4 |���d��=�y���%KB�p�rbK�yD`-p ŵ]�I��@?^��;vr{�H��²���Gkݶy�-�ԚC����gX�<d��۰v����p���X�])��C=�ռ~��6��Éذ-�wؿ��ڒ'���	�] ğ�̓�	u�g��-8hC�����+�H{/�S���Byaܓ(�B:���q*������<��7[��}�å��,�$��'��A�%����Z$o0�[�n�|E���<S�x,xb ��'��Sa�X[�5���y��Z��b�ǀ��γ
D���Lև�_����k�1xb�ƛA�I ��0�y&(�_�>�<�1��V�A�q���X�J+�/f5�r
�u� S�R $���� ֕����K1�wAP�+���V������4�����M|�YgZqh����n�`�};]3�=��}�zy�9N��6���6}�LO��oL:\�f�lϱd�j���)�Z�{SV����֘�Ա%1]Sub`!���+K�-�,�$A��l�q�g�U9a�8�����3�N9�6s��I-Z�9ߛ$X���]i��9�L��� TG(:=�|/�1��c��5�H��4�F��X�-Pӂ�~Ah��&-�V`�0��5��Jck|T\_QJ������#M<�}bMZ=~e�s�6z��^��K�Z!v;�hT$�֐Rc��<�^��敟��@9��)jH�C|s���ח/G�+%{:��x���8�=�7e��;�s�\����?�{$��p~���/�L;�&M����t&�͈z�	�{y�x]�oQd�?�B!�!<�)T�$V�4�u�<���%�v2I�"ǖ� �#k���Z�|vu�����g�w���74����h�6�_s3j��OU��i�!Ty��uV��qG��	-�����v�g?,��Q �w�7���s��cmN�/KC�F ��,J 8�2����%bm/�$F2y�1�Ij��D;�D���p��]}-#Y-<���B����I���S��4�=�UP�B0�!k[m	�T�:귣���+��w ��� �t,e/���;�Xo�7$r��wYd�����w�q�\�g�6�Xu�O�g��?����Li7V#}����֑�oϚ/-�U=т��"�R����rŲ��l��e;�Dh��YB��aa7)B̑�]މ1�
e�Uԑs�N�_�ּ�0��lG�[n$l�P��;r!����CuR���X.��a��V~��X�o]�!h�>95����7&o޼s��Shf�8�7*�*��v����,&Q�>ͦ�?����c���wo�Q/�&-J=�x��ħs��?QA�P�֢��(��ck MK�]G�[�}�����^���zҤ�;O�2�}M���K�$�s��]*$��*5�ԛ���n��;���@����_Q�� B���o�ݣ|h������������A�A��AV)돜2K�l~��_y�!�{��_�E�PD��d%��q�����T����	��Z�W��Z�����%�fRV���9��V�f%�}���Ý�MI�0GP�t�J���aI瘮��m��J��+E,Vd�/�r(Um�DҜs�Qv�s����&L���*p�|�
[�jm��9���wtUUh�ߦ�[:������zgʪ��o���E6��s|B���r专�R�y�Q������M�;�(F�W6�w�i_|��� n��f/�,���B���&Y
�}L�H;�ƌ���v�V��"���.��G��o�L�*$H%��]�P7)������J���4�%#� Bat�g"ڧ�;P�3�$��'���_���l"Q���44�v ��ݾ��o{���.��rX�4���_^_G�]w���34a\��^�'����?�����ČG����g����̥qݱ��B���̕j=i����[BC~�u͘q�W��;�8�y�t�|����{����k��ҥ���w��a����;���g��i�r�j�Z�>c�{oY����u����-4������P�L>lj�ܜԩ�_-��n�L�^��/8ߦL�T�����n%�~�͆d-Kel��^��^���1@S�����\k#&�l?��O�/x�oR����ы�Q�)iӇv�&;�H&c�s������Lp��( P.1>�`�w��OL�	���X3���{�񓟺P�v)�E�.�&1�M{!5���a*���E�A} (����J���??h�q�>�nD%��CH�������3n��F�S�r l`U��J(X	���Z�b$���7�#X�?J�����|��|�7����b]q��y���BG�&�\l5ǁ���������e>��H�ճ�/^�:[��'ͣ�"X�V,��Cfx��'�Xj�/�D�\G�	�'	�#����V��Y|�^B6oC��v޼��k_{�M��e�tնm�l+V,�%�?b��l�,����c'�x�}�s���ȍ�SA������/4 �۩�����}����Q��+��K�,�ו���
HY,&z�"@�8P'�W�d%����v�F�l^�W� �>��j�/0�3���[ns�U��w,�Z@���)��wн���)�����[֯��3|G#X��<�ǀ?7E�����}>��	�#�i�A) ���0(�} o�h�����6�( (%� ��J,�������}3YN#�5�w���Oh�.���_�}�dK9����U=|QT�O�-t>���4����VX/eֻ�y��m[69��!3���͵l.o��Xg�{j�*/'�z��?�h���j.��_��?
=�����3h,@*xN��f����J�1}�UJ}�}�f{����򧞰����iV�x��!���?��<{� 6����
C��_�����|�+�G#$=�]W\�<-ş����E��i�b�̵`�7�E�l�V�C�����_��o%)�`���i��Q�	�"�~l�[n���q�u�G���FZjD�#m�����?vFslɆX����G��\�5�wu.c�Ӵ@F ��W�(� ������d^o��G�G�W�.���_K�g���w�!����*Ҁ?��I�0N����D���O+��{���"�u��g�������÷���>�N�G9 ��Cq���g��H^c=#�����g}#�K�?�7�\�Ry�{�a��{�9�Dp��6�?ds�e�}�͞��x�G1��n��P
����9���M�r�8��T_�k���۲��-y�!{��-��zQ|fY�e�lgϠ���q'�j��z8ߗ��e�p��{�s����I�OU@z���	ƥ�H״-�F����"t ��5�q 	��f�NL-5�rů��*���B�i� ɢ�;��{�}�����K.�gD�yN��IS�ZV�,�}�9`�{�+���gV�Z�w~��c���9����p��O'1�D��{����h����5�s��� a��������s�T��5��;�cF��so9|��C���D(?�e8yk�>��p)#�1�ozӛ\������[xXq`��z%k���\���sө�elȖ.{̖=������i塢w��첁����؉'�f��y�z�,�,��f_3���4�����k�N�6Bg>o���]��c��T�h����6uY{�l��^��R�����l��-60h�ik�����y�?&�g?��kq��1� L�/~��&4ϸ�7���dS+$NL� ��9�|�T����88���� ��^롃q$�H�B�����1@?|4e�#�U�(���h	!m��8��m���?��'��GGçp��>����zVǩ���G5�YNz�/s����8��P GB�n lE}iޕ��#Q5�&c�H2��(tX�c��q�OE�R#�۽d��u�gl'5��u��CNH ~rB-L�o��?����������h*X�>�j��p�c@����f������8�k+�z��%��ښU+Bu�rj>7�֮�d�}CV���-o}�<m�<���d?���u!+ 큫����U\�3�����:<�䆯~���O�\�+��_dCfҝ6�_�IJن�v��'{�*@ʅ	_�0A6����*@,�0A�C[ToV6&�P�D���׼�����PWg�h��.\���V[�xbU��u�<1M�E��_�!��K������V���p�bR�$9���x'�h�h���sEg���
e�. �xʿ��}���.��r�_EH�Sf�d�i����u���h����^q�hȝ�P4}r}��a�vCͲu� ��m�\��5s��w|0�l�ga�`�C��/ Jڗ��%�A�p~����ۻ�CgL�I�'چuk�FQ�u��r�f+W��J5c��vۙg�k�{����k�-]��n���m�������T�s��q��?�c��Q�~۸a����;l޼S,�.���Ox�_b�k����m��V�u����l�	��#���&���|����	11�x �-�_����:�JQ�Y� �Z���(K0Q4\0@����<M�@��qBSi`������Y�ȝ�q���]}/��������D�ƅ�u��1�{�IJ������<��T�����d�ǚ�(A���c?.���j�����Bz1�-KNV�֔�Y���؃�����E����$vՂ �4�g�c���aܘ+�p� ��ĺO|���u��,p��"�/���l�#��_��N9�h�1�[�أ60��� |��@��u�u{�uvM�_�q�wM�����ƛlŊUu�����p��3�������o���>Գ�毥v�s�t �Z�V�z�~������n�T�֭_i�}=I�D��-ڪ�i�m�/�`'�r���M6�wh�C>�4z�^ >��?�&'�mTB�LR0L��E�z���d����q8����Z��Z����+�tx>�Ef2���P�lFۇ�G�W)�v`?ҳ ��>�J5ǆ��y���P|�`��)���� 4�틠m)�E�)	7Y��W��9�k�B��6�Iܞ����z�XP�^��i�~��n��KV��^�*[�x��k�c_@���o�i�J��;o���8�>x��Z�<�zz�0 e�=���Ga�v�����~β�N����o�b�r�	Qy}Y����?_ڬCg�'?�1+�,m%��o�h���ݶy�:��� S-c=�A[�j���Y۸��iej��ѫ�O�����L� q��lp���7;��������ϙ��)�ub�w��A|���3�n�k9RZb+��H�w,_zH1�#l�/>#�p|�a��d
)������s�|�|4�ǳ���c�Ɖ^��k�ɇ}�u@���k�|��������5����N��`lEi�]�u�N��'�G��6y�Tۺ�ە�U+V���	l��������w����1k������i�{���}�v�
+��i�N�mg^��v��m��m��ګ_�jN4    IDAT�z��=����N����F��w^�.����)ޜ�"
ɹ���8��e[���L��4g�� J:�xB�	x���?BVj>��Ku�#�>�x�!�G�/*N91����N���������=�C�8�g�b�;��{�#f�Y�kV�p �8���oK�\a����M������ezh���k��j�=����G��V��τN;h��v��U�Cֳc�mߺ��wo�Ri����%ˤ��/tÆͶb�FK�&�;�����~��1�h�$[a
����O,�,e������׻U��H��J�#�x\��}�
b���8rM� I��~��	��磈'ێ�!
��V|SK��n�������ڱ�{L����C�N��X���O�Mq�*CQX(~�;{�R����l˦��ݽ������}#,c]�{G�=��%ֳ��.���6k�l�T�v�O~j?��-����)��%cx�:|���QU�t-ms�εw�������[��=��a+�l�L�f���@����c�©6�9�8@������$ƟJ���DD�"5֮_��f��0��deӡ��H����?�m=~�31�p��V�+ �Xxj�  T(Q�s׭�����G�3!���c�1�X��V�]��ʏ}���O}ʁ���\'J��N�qQ���8�@	�_�q�h�V-�e˞t-ʇ��\�_���`�N:�t�{�)��uX���]��=� \j% �8�VU=�VO6D�,���)S�S����V��k�����k˗=�WS�5a��z�iv�9���鳼�@Ov%�J���D�/Z	�-���� ��N�V����J-s���7�5d�9�q��X�l�+�EV �1�OTq(t��1M�HłA����9���,h��<�x �XޓwW4�"|ؓ���<��x�c#G0>u{� }@��˟gR4?��=^t��T��Ѐ=��v����+�[�J^HH�<a��v�ة���5���<��gw�ү����s`W�lQ�_]��JE��5�bG�������Yg�n�Ҡ�je*؎�[��[��'|�t�T�e;�X���y�ų�0�lU�'��/�ω'���]D�ȩ�yh0,.�>o�1���h�fe�h���]���3kmK����=���TB��b�e��T�#�u���Z!����eK��iU��ݳ����Z�]�I8�	�&��g�P��������,E��	=����ՙ��ނu��ڵ���c��>X3gf�"��t�._f����~ *��Ƚ�g��o��Uw���(�J}��|_����/8ߛ,PB�hRJ�ԩVC��޾�����=U�/����W_�@�ǂ���+}�X����_yHQ
,���ĉ.��9�� �������0�S�-�]�z�gvS���P�b�W�H��0�U-�N۱�k�$B�<���z��р|�cT�	P�ު�p����+��Q��`�<��Hй��P�^������_w�[t,+��~����o�B��G}ܾ���Y���^5�\�~?�����
݅KGN�ҿ1��o�P+�F�&L�I}��W;mCyg>��eaB�l޼ս�j������1hj�v���A$;�ݮ����¦�|���f�����u��E/��pdƺ)Z� r�YH�m���RI�K~��a3C�ocl��Iy�V4��s�єw`̈��Z�ot�kG��hL�	5T�ߎ���l�ќo*9��7~/@�3�UnC�[��O�c��*˺1���F�&�4@�������Y:������<P"�s��@V*�uMԏ*�����^U�U����Ο��:"��G��t\��ڱ`b/S��w��l ��_Ia��vK�N^ټ���!�ε��&{73U�,�"���3"���==Ng��O�������3�?�{U�er�w ��9�|SQv�֊ ��kA�����z�^p�c��G�'�hB=�N \i��$���MD��JU�z�J�1h?�z���ΧV�C���0S%yQ�ᐩ�F��5K�P��| ��H���I-s6�j��o�AJ9��y�X9�v���PVl�Vr�	���v�h�}�{�kK�� 9�5*�9(*I���<�ϕ �2ʄf?�0�}�o��"⪣�KZ�?� ��GQ�\����C�k:�=y�s	�x���8Fu���
#�{���zdN��\=�����I'�uE��1.���}^��н3��gýR�`!��F�w;����߬\����!�������`;�Yw8�� R�l*d䖂êqQ�����'���� e`)���O~�K1P��k0���Ь�Z����uY������/��K<;��z���$�8r��w�'�2��1�uI��nu�������f;��X*!R��#�*!�ZD��9����ƒ{��۝��R�S_'I��:�\IJøގk�{��%PdQ�Y���M}�����E7V�˳���R*����7�(��8�X���r�����%y�w�q��ؒ�] ��v��|�a�8�9����&�KR���_ʹ`���Ă�n��(���;��2�j(՜��10��hh�����©q�aځ%1��W:�����& ,��iQG�k�$��(
M��.����n�4��q-� ����S�3Lnh�^L� %�<cA�CM��%%,Ne3rV	��B*Z�#-���H���i�����4��y󭷸�[%k%�)M��c���;���Jƀ��&�*�;�I<��6�~�r�&�����+n��F��I��=�w�y� �`Zq���)�����gkw�-��땠Z�$9�S���Ny �͟�J��/>88�'�h�=�H߫���Uq,悬b�Q��P'~R������:��4*�uKh'-i�T�d/�I���z�p��`�9t���c����[�a����:|��)�<�n�jA�G�
�t��b4�J�ĭ�r�w&NG/��D�o��w�Q�4p�	��4B)8~B�`�?=}��\RW��O���P�v��1�ƢVm�F�_�E
��@ʂ�7l,0�	��ӤƋ�Ն�����8|���t�Q?5~D[�n���$� -���/�_�\��o�y�V�֧�㿧�6�S\��)�d,��1��3>�C��D���1�ז����+�Hc0�wP䞔Q<�p#t>�񏏘������j�!���ZA$��t�M'�%����.��{/&��?��S4vj��9�ƨ~��0��̹j%r �p��TI���F팉Ŝ��o,s���v�]�a3�q��D#�����y�E���c�G�̹^��_���GE� mC�&	o��%���9|o��mN��;�GμUO�}|���ռ�, 61�<
�y�ERu�&}�1	�?Pn�~ 5�6�Nh !�^c���7���X0�bJ�k��%81VXI��sٝ���c��Z��<vXJ��6�ؖ���5��s-���}ޑ�Wt��>��{����M=���s	����#���[*%��L><Y�h�`����j�P�8(��c�lοE��k����HӚ��L#�j��PfA� �Cㅴεهs�h8��f���3�T�.�A6h�Ī��x�K_��_o��ݛ|���}ڙ�.���K(�H��_�����YG��ӈ7'�}�[�����Z�%�j����p��&��r��`����(��7�_�`ų���ʺֆ\H��Y��]Ig�� σ��:�hr�]�!a˽dep�7��u�[k�v�DϠL�՜�=���/���Z�7���/ņ[�ַ�o�(�MhY�g\v��۽����u|/�E ��Ou���]4
3)ij(q����^�B8y��� �]���B�'��F�g}�}�$�V��6(��������J9h"����kv.�E�*b3O� � Z���j*���U��lp	��h���z�����k�'�3s}@�{�N��h
�-	gv�Ӝ��J�½�������v��L�,��rSI��	-z�	��d�k�	,�m�=�>����
��y�K-�f��ˢE�p����ޚcͫ�|���3��:�_|�cu
E���<�p}���{�ܘ�z�K]KN/�����|
l5�;�m�Gćs��#k(���k� 5�w���5ͳ�}�� �@D�����}���,��U��4r����a�N�c�}��Ĺl	�f���]g�aV��%���ש� Z�j�qԹ,�봇4�X��$���ڔ�`k3K[��N	��G�^���":���7��ɤsP;�m�X̭>��X>ZԊr�i�+C�N��X�m�ϭ1ֳ�����Ƈ�cݐ�G�a�k���W�q>
oe^Y7$���_ �O�'��ց�ќ���F{���H�VS:᮫� �(d�1�K���G���{�ð��OJ�H�5d�"n߮��j�����5(�_ᥚ{Y$z.�����)+V�\:��[�:��0aP�p��q�R���bZi����Z�UfN���ŋ��5�I��z\��n8\(�Z�f3!<m?PA�
�d�<p1o�9d�2�����[2��P|���^��/ ���r���AlA��'`�l�*D��e��iNc`޳��c�T>��9d:k|��~��e����{�U�k:�~K�.��2������C���x:LUX��|��zA�v�/���g�9����E��e#ϥ������+�|߯��u�^X�-���W8�j!J��s�,)*��%�yX#t��3d�Ha�<�Zk�fَP�'��Tj�vM?X��/���l` 亠t��������fQ'�_�iH��gsA{��ET*A���	�삏/�dtuM���m�G�X��Y��5�"r$)����`���18�`k�O����o�������c˪����6
���v�?��ey0/ZC�B(���ؕ@˩����X��<�@D��Ɖ碥���|����xʊ�T8��=��كs�!��}+�_o-�.�ZPb�v�':_�[��["�CG������mw���g�a�C�JV�r�k�o�	C·"ɔ�r�c���OP:�Y�Dw��f�h,;�����eѢ�5��[��2�vH�pS*���<ҙH��#����zz��9��*k��2��7W�?G����i�P���c#$X���A9�c�kԲ��Z��z��3vJL_qSi����3n� V�\4�.n�'�I{$��a��r���D	<	t�ݓ�.}�.�5XG_�����+ϱ>{੓���[N�Ш=|����,���-T I�5�kX�D�L	����eB*�sR��E+A�č�[�#�	в���i5t�#�PX~ �O�?�"��-ʸ��Q
�|H|?�2�}*�O�4�'�@`��P�	��3�-4��#�wIݓ�u���{����I�ä��j����+��+_��L�4w8IY�h�ī��� E P�����P�Z�5H����t�Ӥ{���6w;�2Vڧ�{����힯����^f�45�9"����ii)7ɉx��7�R`�M��m6o�E�p} �� W��}^J�gQ�I4j�l�r���+�%A�t��(����^���{��QC�lҫ@'as׸��e�r{�q�^lq��aD�o��*�u��-<�,�o�%�޵�M�4��e�E�S�vJ���B�ּ�1��=���g̜����{�N^0<�=�Č�8a�k�z��k�>}�o.����pg"���r�
���d3�������S$'}�{�sm�c�S)��G13�Ac�yGF�D��]�����H�c�v�>���>#	����{����Ώ��;�M���T�t~�����Tkgo�"�ⵡȣ|�^AR�	?Q(�$�Y���a,c[n�3��ц+f�|�.�G�A��E����vy8���o�����w� ��h5�/zE��
��=Ĺ�o�g��	����,a���7��N�����3��a0��7�a}�\,��_����w�s�K֟�w����s`g�.���B��f�?���W��Ͽ���/�x|_�I�>�>��p#�-]�G}ԋ�!��X��$/!����!d�&�DkPן��4|�\���`m�FN�QP�u����p�÷Q���tO�c�v�����������d�b�1�lf=�z�{��^=�}��6����@��8�����J���k�j?Q���U��N�8-����9RO��:���^��:�SW(v�c�˾dL��ȇ�ͬX���	����n���d_��?��{�'��"�:�'|ods6y�A�y�6�ݸy�w�A��r��B#���m���5c�R��l޼y6�E^�&��o�f�
Ϛ���O:�4;��6g���2����#���7��<>���C���?����?���Ԑ4 ����E�&QO K��'5�ݱƺ�������C�'-p_ܿ�5�PX+hb�����x�����$�v�s4��2�&`"��}�)?��=V�����}/�Cs�s2Vʒvn��|
�#<�2�I(u��'��4y�Y?��T�z[�:�X�`1P�ΡW�%랂����~�m�C��W�%σ0�3��/���z��1����_�Z;���B����mt��rQ�4�����$�;\��Kig��8��3���[�F�$��Ϝ9�.y��v�)'Y�4h=;�ۃ������>!D��P�{�̙��9�γO<�r���o��v�Oux�I%J���ϸ��`��ٞHu�M7�BQ8� B`o�v��@��g�T�)vp>s���TH�Q����k��ۃ*2{�;�a'�=ޣ[{{lӆ5V跮���xJ�V���� �P7%���s���I���ȭ�
�쩕��uBI �	��s+�K|=���uS�����\P����~����Q�KKz(����g�A4��fO<�����_ن���EG�;����K_�J;�i�����3�����X�Ԟ|Mn5%�I�����=2gh�^���eo~����X�V����Gy �Х,mIĠÎ�ݶs�l�}�)�����d|�_p+�L�^ij�	��B@K 9�@	"\G�9ƪ9�������h����}������ڶ?%�N��J�^�nmw��|���:f|x^�8�qکf����{mӺ56�W0��)�x�\y��@瓊VLuج������X:�a�6o��v�=��ɤRR'��w�e�)���UI/|+�X�m�v����*��d[�s���N���?�K��m��'l��mǎm�ˇ���ض�������/p�'yq����5o ;�������G����f�?!��\Ʈ��]v�	�[�<d��M��a=�M�a#NU���P�6o�j�r�zz����y�{��o��>�
�BCIJ�FS�o���1�X�,�}�����4�i\��7C=�=�Cy��}"��Ya9��Z����[��P�m^�����[6U�t��QT~<�<4)��>ڮ��N�YGk��l�|�mܴվr�W폏>�+�N8ޅ�nr�%j���|�9�9���|��������+}��"��p��|�	�ʨ8�g}=�m���l˖��}�V+���O~�P�f����[�k��v���d�Ϛ�>GJ�C5������1��/�����U���#f٧?�I+ؤ�v����K_�+�ؚ�O�P1�Ϥ����o�W���!�������h�+W�ts�E�v�$oȞ�/QB����x!��(7I�g� P̡j(5���������)��=j
:P$k�}�{��u��V+Z�<`�6���m�,[��UܑN�r�g5�\��8�	�TƊ�)v�Q�ڄ�S,��t���7ڣ�?|4%v�ǘ��2�����g�����'?���wB�����>g���o��(~D"  �t�l���;��C��	9[�f�����~����mɓ+��s�-}r���%�_��I�z��-[���4�.92��`Ⴏw
ok�1�s�e������%۶}������i�t�֮{���{��e�����    IDAT�b�o�������csO8���	��/���o�' Iߑ��kV{$�LH�\�7�����G��J�ߛw���G@�}��Lo�P}6Γ�3��Ph�r;��ӬZ�L�d[֯���sT���x!!���:���9G[��If�[�q�]�MN��5�p��c3�PO%g�X[�k��N�o��o��ˇc��K5�T"�pN�İ[���_���v�I���i�l��%68je��R���\j��D�)XG���G>�e�=�._���ڨh$��f̜��3���7�oo��cY�l�a��UW}�2���Y��������ϰt�h+V>i��`����m���f�&K�'ز�[�O�+�����p�0���D�Ш�Xl��p-8@��r ���`e	s��8���z����N�V�K�z����1���Ͼ`ݣ��š�rѶ�_i;�n�|�h��̥�g=�W�x�������?�c�z�6a�:�_����ǖZ&��������/'� ]�^�erxN�{��]����T��}��\�(�|���=���7?��O?ΦM;Ȟ\����RC�\IY���Ǘ��J��ne�Q���������W��ei�z��
0�q�o���P��c���|�*������n��[���e��N��i�2����W�uk�8�j�v;�Գ|1�0�pH�R"���p�͋�uHn�{��_zM� ��Xi	q�X7����f�����5(�u�����1߯��S-�\�߲v���������<�����pNJ����MʩSژ�+�.;�����I9�a�6�{�I�>{����w)ɐDټ�U��K/y}=�����Ɗ'�+�6��|���n�Gp�Z��~����I'e3���_,FLeϜ��Wm����M�ի��f���_J���E��v�?s���,^����1hޅdls��9�=퓵��{���Gl�d��J���l��2��l����D��Sy��9`�W������ۼ�^��=1�E�VOU�X�Q���5k��0��;��]w��G�@ H�h�1~�����2�u����kd��x&�M[�0k^e���f���_.Yy��6�[e��[-�*:���s�?r��-D�0\2m�s��	��t6���W��	���h5�8zF���ڹ��m��]ٓƯ��4���>X���Ϗ|�#^�{�f{�ޟ�ԩ6m�[�&��j�O����-yb��Kۺ��N9�l{�%o�l��Ճ[�n��>�4���E��,DԠA��Mo�y�βJy�V>��OD��MV*S�+0qZ���wز�k�З���>��?�~*�+�-�_ř ~������淿e+V�p�W�Iu}�Q$������ZV�B��~�8�$�U�V�+ئ묷��&�3��]��fB�$J?�Pޡ��Z13�fqdh&di���o�����%K<)ʅ_�#@�Q(�(�W�J�ñ?�[��Ź������bG�9m5��F���gj�fգֻs����PiЊ��z��T���A{b�S�}G�]~����G[�����.[t�b����w8���uj��L�,X�B��n,��90�9�ܳ��^�5��|�=����z�2��-���UB�g&�����)���'�EA��?��?{B��_u>N?�tC`Q@��G> I:J�V���D�rm�6>��`��M��@M���ζro��};mݺ5�ӽ���L(�P){�j)�����[��pJ�lαϵ�3�r�fk׬�k���_�[�t���bv�m��b��GV/����|x��.��"O�BK��Q��i��fW\q���u[G�h+�z���1��3��8M^x���6ڑGg��=զr�z������
�Й�f+���)��Ќ�'kNN �-o~��ܼi��rY{쑇��?�gO=�ܵ
�M�2ɘ�SO9�;�X�0�5��~����U�a��kQ��E/z�O>���'�}�l��yZr�&ܳrW�?���bT�=���-��sfϱt��e��n�s��8��R&�v�5ۤ�����̆�;x�t���ٯ}��v����Kg3^<n,���Rv�BV�s�ᇻ�O�{��6n��A������ܕ<W�pL)���~�I��mp�����>۰a��{P�3���Km�aG��I[:�����{��7%� ���?}��?? ��/X�`qw���f௸{�e�v�An��>���b�y�F۸q�k�8c �9�g۔��Z���Jռ�%}�"����,t9�X8,~QM��n�A	 -�����Q���C�G`�G@>	��؇h��K�������i���JRO�`;��7�{�dC� ��syotB��2Q.y,�P^Y �[��f/��#�K}�TЯ�kO��
@�Wƾ�J���[.���'٤�]6��ok֭��[6Y�@�G;utu�o����������sg��46l�d]��R�|���h�\CA&�:�d�⬁�g�,jF�Y���-W�w�������ކ��rI�Z�B�������� �-��1�ݻǘ3~�d�� �>�F8�N�T��x~��E���?OS~� ���b3�\����/��k륤�m��nr�q��#y@�=��I�1��:�����_o(٠�`a�D!,:)�X�0V8f����^!����S�W��6�Z�����Qb�4y�$��N=��<�v&v��8�H�K9�t���v�]��D-R�	��#mGf��'���\n��Vw��!��}����kk����
�=K���c���n��ִ�Ls]V��U-nըf.O�2��}��| ��<��$d�f|o��q�!��)��B�k���.�GA��=��c}c��@_g�	�N������>˻{�96i�D�˱��W�xwa�=��?�w�����������颜�E��¥M����E��rJ=`�Qga@�I'�d�6+D��.e�n�:{rٓ�uTke?��^����|���������Iǜ�$���/}�^�{�g�������Ox�F�9�:�Gh݇it�x6g>��TÊgv�(�\:X��%}�^a�����pކ���z�*�M��aһ���b�Ja�h�T椌QK�ݶ���H��[n���<x(�SԮe��1Ӟw�q�QC���ֺ����I��� ��Z2��g����i��l���-�wh�B�K,��*�)$ӏl���W�&Y�.���+�K�I}�At!�$�aʱxT/����Z�*?�7���l���z��T���(?�o�G���V�F:sU)��M��Ϯ�<�(����@��Thv��tٓ���t���l�T�Mq�q����.��K�ѽ���5�y�G��H>�},���>V�s�\.o�	���A�� 4h3h����i�jq����=P��Z:|ہԮK��z�g6U�V�d�0� h�w�����/�ܣ}p�7 �_i�m��6����ydA�:_�$��03�}g��3�v���iQw��=I�zvvҌCᇲ�d;�c��c͓�"q"���n~������s�]H ����[�s��J�(t����9��\�<��Q�~���Iڵ��8nMg��Ww�ۃ P���H����8�"N<k��W�pfL��������t�v+��N�'�^h�� ��&�|�6�I�Rr����gqxƐ���
�5{�Z� ���\(t_Ҍ�i�hw�4�H�HׂD�F8�QC&#�i�${�(Xh�p��?�� Q�8mt9��=��,�F�R`���H��I{�������ꫪY9�Te3N}%�qR��"����ZXm ��3�;�Y�A�|b*�N4�D(Ś����8b%^+í��÷��0�`�?���`j�T�H��r+�|>�A3ޟ���1���F��q���u�b�|��i�E���@0r�E�m$�4�a]�8Gxb�oT6C�]��� ���[
݅�5�Ȭ�al0����ݵ�P�C��&l܀lB�b��y� H�ูs��_����G� ��|����ځ7k'��c�s4�����"��H���6����|�p�5J���F4��Q	u��Fo��s.s&
A׌��Aɛ	��g���]@0))�b ` 2����
�9K~�z�9=����]�曗@������/З(��I�S�%
�5��`sW���� ܓ�I�fb	Z=�����@���v�q�Ջ�)��y���k��U[�8�!�����hB� ��ڰ�$4^��a��*��:̀?~�x�Ŗ � ����b���;��š�qmX����M.����7��4���f�Цiw��o�}sd��j�Q������
i�~�H#��$:�g?��Gy��G�^"�D�i�wը?잼a;���w���e/�g!_I��Hӗ��"�#����<)%Nt�~��H���zaTJ��y�4�yXL�7n��S)XJ�ЇW�SFN-�^EK�okĺ�?�,�?��<h)��g�����������w A�5�@2v�{�����o���/�0��X��'�ä�$d��7"rX�h�Тb��Do5�rI�m#!�nc����O�n�d~�k��'y�]v��#�S����6��V~g�5�׽��노诊3��)ϭ�h�Q	�=��9</�Bx
��1S?��K.q ��C�(nY<�֦�T�?�C���~�v�d����� �IɆ䨘�ј��\���`l�I�fi��.�b�^`� Ƣpȕ�В5m�����beLc������0eLe0�g��Ɋњt��,��c�. | �u���8�9o�[���mh�с�������<�MT&�DX�p�C�x���x�Bk�)�����8�+�h�l��*i�!��NDD&�z�}����uɌ���{�J���ҾΫ��"(ش*�G�Y1���ַz��O��]�W`�����2�5XK��r������}�c@V)���F��H0��#Ǣ4} ��������=w�W�����Dah/����� �m;��Ԧ������O��ݿ�m�C��<�( ͵�K��i`}�=��z���X��t`�f�i$�W)_	�0t)��`ķ���8��bǵs����G��kk��%��1	!�D��eq�~� �`���h	���e4�M8���&�o|�;��m5L��Ip�o��q��(�y��۳�c�����$+�ͩ�
�CV�Ýު��/j.Q�Ma�d�V8����g+A�O������$�(,Z
�9Gq墴(6ȹ|�(�z�?���τE�j�b��-�,}�CH'�a�/8�����]�v��X�$�R�4��ź��[5�J2�+��#h_+Z,�V1��E�P�%��1pBkС=�C�sW�u'n�^
�<��$�HB���{��>M�R���Q�X�������^�W,�i����6|aW*aMS-����r�4�7���A,�4��c�\s�5u��V-$�<�?��@S���Vϱ��٘�?�,�GqB�G�d��%4��[h�1u�9n��G�ٷ�v�����_����Ų t�	�(�9�:�/�_>Ɓ�~��փ�����pD����빗Ʈ�4���@K��%��"��=�&9!�z�g���0Q���[o[;	����FzW������*9���`Q��^ba*�w�Iiq�I��	��  ��
H�s�o8����U��g��[-�z�q�V^�_�G1!Lrp&��X,{�	���PC��s��`��g��!�h��ڀ7�i;N]����5r˼����'��x�R��OPS����$υ���UO9���M�vϾ���%�{wzI]4���6&sR.���&��8i�Gċ4�Gy�#4H�{����2̳��4ƌ=��C��/}���������;�0w6�p�����w(,E��x��~|��O���1�� bE��p8�'��P@x'~g=b!���3���|���e;�Ph���)�(;�	�q$�F�_L�2�ڇ��~��J��E�J�c�j�;�9�5�����go����6���˓!\�s"Z����!<�����۔t&Ҋ�r�'"FJ�PցZ>C�%Ky"FH� ���&�����L�R�Y4L;͢FHk�f�x�21�)���SO�%�i���������/: �>�E�
`����6I�wؗߏ�1���	E�0?�6m�wN�]xw
�Q�	�j ��Z][��\@IQG
���s����������w��T<�a�5G=V���U�6�d<��z?E��"��(�����d��iR���Md��L�X 9���=���Xʖnų�7�F�  �<Y�R��(Q��bv}�Iu�l�f�:��BL���'����o�g�e�j5/���nj|@��k.�vO��&-.��Ҩj� ɏ�3�K1�9&d�i;�?�6W� k�5��/X
C#BD=V�XQ)--J�G~i.֕�;@qJh���Q@��&����m���x��Jh|d%p<�+�z#��kd�����w�6w��	�JCܟ�'���?��d]�����|�󰁪0K�ħA�1Q��X�_@��KE1�5[�����+SV�q�s�����$�+P��8���z&t�_U69�DU�a�Y��,+1�z6����`A��C(���<�1Yj��O��u��'�d�7���}VhKz����P�֮]��@��t��%���'�����5��o
=�5���i	�_u���PaS)��c�����;;;|a �;�&�@ ��O}�S����|w���b�V%�BT�P�0єp��PBVB+�'II���Ɛ��p*�P���'@�;�/Ĵ�H���Q��9�Je�����@,����yVE^�&y6Y~Ҋc�E`]�I4W��8=UW�x����@�gx뾚�v�'ZNjY�. �!�MTǒ3��;�·R�>����{��)Q]�J�:���	?D{��V,���yq�c˹����c�'�k^=�GN=h�K�^��z>�jmE��AQ!/��$�9�Ƹ؆�@�?p{�.\��B����?]S���>�>t�,��9ȗJ�t*�<hK��o����cB1�f�~�kV,g-�MIF/�a����;�vXDT�r�Lf���|:�쳝n�)�8	�j����P)8Y耇��:�
�m�}�}+���%s�<� R�x%�(>����Gs]=�"������tc���6lp��:{�E+��*���=���q'�^�0)p�gfM���;�Qk�[`C�a�H���`1T��o�����$��������;�$K
��X��O�AEO|K��z�~����y�B�}	ʕ�=���x��9a�u��N���s����~��۶�p��k���7
=�l��Z�ڏ9�h���WY��édS�`۶l�%K���֯[W�+���	�og�=Ϟs�qf�഑FF	g&P ?^��� ��b�U&??L_��|��\�S%P��]W��fϱ*���<�Ѱ1���}wa�h��� پ8���Kt�������AQ�SY2�c-V���~��� �.�v7cރ�NxQ]{��㋢Ě�'A���)�/F��ͧ?��\P��}R�.�)'i;�G�]T�:��3�K�����T�Q�W��(�/�fmA�~������;v�w�̛7�#���k/��^z���O^lV�X&]�'�\b�V���Զwo��`����{��v�igء�fCŲA��w�u���e���.���Pxw3�VC�c�:ʮ|߻�R�l�҂%[�~����{<�'�	�#^,��P���*6�������rV�~�eJ��� Ŏ?�|(�a���.�Q���h�8�����Ƅ;��,�����Ak��׿�NQ�nc��o��h�_c�@��;�ck�x�V�_�-�-V������>h�$�)}op�Ҁ�����:'%p@\8��'�Ē��西�ۿUVk���4x9dꣵ�e��4*ψ����x�b����ݲ�#��+�^�w�(B����A䟀�j��Wi s��W;ː��l������ۭT���N�J�N����vX��������3gz�2�/}�Z�0��8�7�\�](�yS�'ڬ�=�������:�+���G�\�f[6��m۶��Ѐ���&��d�;z�ڂd    IDAT��3`���]����ɇ�����!M�@&��w��Zil���\��_���9�D�Q�5
�=tl� #4�$q���}Ќ�Iʂ�F�_ ���}����[�h7���z?�񖦪��
9m�c�pH8�.ມ}�M�7�_�'
��E�ٗ���z�s;p��g��1s�L����.�3}b_M;k�s��wQ/�۟�2�4j|"������]���wgw�}�7jU*�? �/�B(�.������3U+�6ԷնlXc+V.��[^�D��l6o����y�����\iO��x?�������:���]��bw���f�_K��G�9�>�����@�M����n��.��� ֮Ya۷o�\��:�]�u�[�n�Y���o��N8Ů��
7�]�Z _� my�ƍ��H�yի^� �{*zB��g����*}��z�ȗ�ǚd��T_ ��
�����w6 �Ɔ��;���X�o��}H����w�+�BY�� T�h��rG]+����D�z�Nq��G?�dAU�P�E��u��FT�	�ڇ��Z��������o�AH�r=�&��g��%�g̘�5���|ͺ#T�dAA��X8c)��	��ՙ�O-�AC#�3FPP#3���07�&NX4&�q����d"b"Q.	J�F�^�`��@7�s1�xM��#q�Q�iA��޻����WOq(��k�jY���t�W_���<��>�rP�x�Y��M�Jc�����׭5~�ayy�ik��wW�o�˫͇��7�1�w�W�A���u�Ŏ-M(�i��H���<d��u�d���_�5eʯb��݂?�燆�������M7�p�|���<������Gc�MC�G��9f7L4Ti6|LPg�Ix�f����QGO�- ?�E����8Ё�<�P54 {��G��ի�Xx��J��^fF
�;�?��?}�o���Z~����[���Y�%��:�d�fu䘳>p���� T�8w�~0J.@�9h"�S���"X�6�M�EO�%
ȋ�"@1q���yꩧl �@u��$��3 ��/�Iu<=�("��RC����0�a'ث.��0����7W��>5f}çf�A�������~����ֽo�����bQ[�ߚ:��-��K��<�Lq���/2ш1�]e�������cL<�l>��cӴe�Ow�+LӖ6��ǟ����yo�f3��/��.���0l*�@J����ۇKI:"`y��[-=|�p3c������8���,m�S���R�A�C�台�.����JM7�dG���k]�G����g&���M�TI!�"�'��-�.�5� _un��<
q�|�X�d���Y� �|����_wQ>�f+�y�ր{��,��^ u��M56����9r�5 �V���QG�6���}�|P�.�$a�zM�ii��-M���%n~>w����kk���^�j���g[�IS&��m�$�����u�Af楗������d=�����<�$����47��`h(j�������ΐ���Ō8� ��N��\s�]t4�ܹs-/�;L�>�Eê��&��c�)�:@P����\௳ v�
�l�����MK��ϢH*��1��m%�FA�����V����hH��	2�~�Q�Z]Z��a�����~��t���C�˳᧒8�X��2y�9�G���;{Z�s4�C��|��]��3G�=���>f�wM{'����6�xȼ������N�HF̜��7Ѳ*Ӵ��zZ�Ye�?��UԖ��)S��/��P���G�0�~t�ikm6}*#�ŏ��i���f��LssS�(��ټ��ԯ�Ĵ�yf]}�w�?��*�}p�(��h��1cl��,����F�0dlD5�Rj�
Tz�i�/ �2�0Ȳ
��eec�0d|�,l
�y���}7�ߵ����Oh��;��Ϻ�R1�}�]̅hy�<X�Z��]@6S�Em�C`��N��@_���&�y�1��c�W��۾� ����Ƽ��-�67��_z�x�P3`@�z�*�mNUl�������۫L$��l�3�c�8�_L�>5�ݕ������?>h��/Z�����s�zZΟl�2���!f�W�f�;oϴ����+�j'�j~Sf������6��Έ9���e��T�e~'�kN�'5��xW�/]��*e(��\bU"��r��)p.���
��B�jN=�T�{饗� ����L�w�cU�?�%��^��N�F���_)��.\h���gk���m�R5�Kɳu��s���=7���+��Wz-s��o��k;v��������%ւR�<���iv��u��0��m:y[{��:&u6���'����]mZ[�滧�iFr����k���^��C�t�a�Ǉ|Amm�}E���LY�5����������ϛ��C�d�;[�����7�3ﾻ�������ܞ����io��ƦN3쀃�q�Oܦ/��Y��<��ݨT2rF���*
c��	E--�=��rnfDO�?�������W���(��{l�Z��(�02
�10 #
��5R�]�$'I����V ��G�=���v?`��;Nl���nO�
	��||,g/�g���b��b?ślX��Gٲ�Q�jAk
2���V�����u+͇~`�;�MUE�54�imQ��xɈY���f���jL��l�����y����r����Wjݱ�/Z�h�=���'?�;3�Ӷ��:�/�O7t�����g>��`ֽ�����?���z��N�
E��Qc̸/kF|�M�b��T����c�*Iכ�'k%�e �/!S��Z�͛2�}��kv����g`������m����ݢ�l��a�_Q�����R��B�?�F~?Z.�>���2(���X��(Y�
����qXQo��,�G��œ��>���Q����I��)�FԨj3x�D���7&�n�Z���_�����^5��wXs��:ZU��|��c��8ҔU��:���j���{MWW�Z���2h�E���w#�?�;=��O"x�3<�\p�~��6SQI5/�.v���&[�a��>��4π�M(L�0����8}6���S�G)�Hq#�p�|�@_���������y���!�s��P�}uV��J�T���ϗk����@���J�
HRTUc^�o	��S��8ܞ��M��U6�/�`S�|jW@}��/��v����Z,0�o2�ԟ����~ �?cٝW�-�L�K��U� P*R�M`�ޢ�T$�B55�S���Y�<� ˥I�$ݓ�l�w�3��N22��0~"}er��*󅹄��ء�m�Y�V�N���$9=�Z!�x��}��+�@�t��d��P晲s�ռ��u��4�4���I���|����oжй7�p�Ut�r�<yW�T�Ϝ��Czx�J:��x|���wW���B!�|�!>������U���o[ϊq�zy��4x��ŋ�Ut�����EA�Sy����T��iXm~��L�l(����k�͙��A8�� nZҲxO?���JQlmb��ֳ��ci۾(�d� o] +��o�l�w�y�n82����¸d�Ӧ�	 �߷��4�8Nm>�	��N�� �%����Lj��	��1Gw��{��ލ��� ��\�YʖM+�W��������)���.��gP(l�p�m�ؼiQ��ś3^��s�̖R��e� �|�?���i�(i�.G
�"< [�3�Ea�1�ָ [���@V�1'F�t�_����A��}��-��J�=�5/R��Q�F�8cE��9��T�=k��>�2{Q���x����I��}��r�`/
��!7_2�Z�Ƚ�KH'�I	�=��y�P��u��9)e>�{)л��@3n�eW���d{y^29dА鵵�w�O�2��Xl�iYi���^r�%i�P���2�u��p�b&GY�dA�B#+��E>���m M�g!N���D�p_���{�9��]ֆ�g����V��:�'VY���o��;����,O&���%o�k��l[��WXA����[o5����=�@�a	o��
�@���)�٤,X'Z:c�1mf��OA-Oϥ6���U�/`�����R����n�=2!0���f������<�J����?� �?�ܒ��u?���+��s<2���;��sm!# i��3�5���� BN~5�����IgO������H����)����d�k�0�k���y�f���4L�N�b-�Ħlz~�Y޶�8�:s�J�3g���@>���yF}�����K?��/�j`
Ɣ��xd���<�U��~;>�	�i��HnZ�<d����u�.>�8��b����2�m(ֵ�N�,~iu*��,"`ON?�}�m,hr�9T�ŕe�=%�,�[\"�c��h6n1�Bl*�q��������m2��ҳO�4�o斲�mO��
�;u
����S�>m��WUT����y��l&)-�k���x��h���r�=�	�]*�g����q����7�^��\��Qq��ѥ�v�`�x��z�H�\����SbN @��w_R�Re�} 2d�,�=�.�(�~���chqrޙg��>7Z�>K\�b�-�1�Ϥ�d���[6����c2��s�O��g��{}{�F)ɪ�QCCq*#@ԩ�J~b����w�� pƃGKJ7��Fź�]�}������C�e
Ƙ3)>�xP d��ٯ(�[/Y���d�Ew�O��(��N6�P��&�_ZWՋ�����4��>�$��92a ���
S�xJ���j�An�� (
E�k�IG�*j�T	cM ���u���J�rS0ڂN"nA�GQ����d|x"<'9�|�R۸�@UHV��R�6������*�Y��&��
�G�bL��8����]�Ck!��뤸v%��'�LjL�����di�&s�����҆��|����7�W<+� ���E7OR}�1�wJpd� �6m���3-��d	���'�p���/Y�ʣWF�֒�g�jf(�M��?8��,���3�z�V�T�2�}O��`��KT{�q�x�������^a_��`�^c�6U��Ŀ�E�fƈh_�oK��simm����)S�b��og�d�Xx-� �u�]Nյ�e�sf�YH�G��ʱT����D\�xg�ϱ�\���?��u��a{k��`|?���|��M���?�����pc��bG/rL���	@]�������������B���y�~ �>�:[�L���}{��~}}�H
R���񂠜Di���������"�2t�;�ȋ���Yw����nv����3�N��q���F@F�*��z(}_YW�||�Z��|?^�&t�,X))�����:�w��7X�^s�g��W�j�	䛗xz�${�1��Dɸq %> ��)) "�^Jo������/E��3�%Ydb�0�k֬�^s X�c.�,���7M5)�[ލp@^�"�H{^�\�EJ�>��-�������ű��)��_���@�)��N.g,�ׂi)3A��I�
�[�wJ�k�
tt��o}%ҁ%��r�c9� �Ud,���J�g��R XԎ��x|��tM�����/ZŢ͐���O���>���
��e�5�@���f���l�o���<3|�a�2���gPX��Z�?�Q��8k���ڂ�9����z�QGٸ��5�*��}tϋ҆:ԚBy�(AY��R�2p�K � |�M��K<��ISK����r�
�?�D�7�H�~�<���=��+�����9k��e}\�'��ε��KE�6��c��갺y�|])��xc�l<�ﴷ��(�[�F:��N����b���g~?����Am?s���a�R4�.nHaK!
oDm2���d e�=�Sy�:s�E�*>�2��X�qj6�( ��L����ܝ8�dIZ,�A��U�h)��7�{��J��od�5�CX ���{ �@��թB.m�*�Y?�ļ���nu8d�w6��!!�6c�!��象� �x"����������,}ι��=����$_���e+�U��`3纲A�lN?�ck�[��c���UJ������������V��D� J�C �~D��PV�A�+D`��3Go�����!N|S�f��D��p�}Cn>�$0��(*�/Y�X��/Xʌ᪟α�*'����d��k��"� ���������s.M+c�k�RgϞ�ND`O�	�-ݚ��d^dy���Y9��h<cP���衇ڸ�G���R%�̢.?�Y���\cEϡl#)���Z���amm�m%�O�����d�?�kd �X��d[ @���� ��ȹ��z:��H�:�`�m(��Q�6֩
L ��+Ț�Z6�F��~b���2b�� d_�m�@�����o�_)����Y	xc��I ������Y�� .:��� i��Rb�����X۠5b�?�я�gB�(
O)�xU�.2$\�����s�A@A2_o��Ft\����͂s<����{sv4��1��O ���� ��/À7��IW՜s��f���|�i^ޡ�͟k�H�C�"�,zf�����]��+Gm�0�JBI
�ˀ�U2��}��naݭ%����_�?V,��SD����
�m�`
�@�2��7����s�)w�7%%e��r�-�2"�!P�����L�����Oa�����?c����k���8�kg���O�1,�Q�F���41"����ǈ@�g��W2�I���\?�D�Ld��Vy�J]���|3>y��_��k�I]�O�N�VLbW���<��kkko):�<e�c�����h�]�0;���Y�JU�u8F\m7G�;�*�{e)�9e��9l�N2��;�;,�s@�Ԁ:Ԅ�����[+?�����9Wm���l��--�������Y��?��mV�G����W�})�".!�������H$}�D�'N�'�W���qO�X�7_�����}�`�h���В{����ߕG)�P�W4����7{��1�}�����̪[�h^с����o�&���O6�w�'PKJ��q�A����L�/ik��A�?�?����4���	 �^�������F��ˣ�>�\q���anPrk 7���	����s 	����K\5��B�?�r.�$�W@� .� �,(�ݦ8�b>�d�'{�TfёPrx-J��	�fƸ�3;�������\�����(�Cr,��Y`C�� ��|Emm��%���h,#,������
*+�$|�ff�*���m"~�}6ΟTO����(`� �7�'=��C���( ���PN��p}��e��{���x��,��Iٜ�����?�NcA2�|i��Q`�!��CB�3$艵��@�9c ނ|)��A�}��'�M�m(EdIVv�\��v�.���)��w.�_��x�����(h+�'S��d���Ʒ�ͮ[TwS�P��g��ם���5bQ��[���& ˆ<���m��
oد���dc 초����-��!(�!Ç��j��T;2������g�W|�8X�>A�6�_�	�����	Z�fX��z
w&�KcA�'���R�$�
���^
��"�f��W�&�C��^�_5��,�w7#&׶앩���Q�x��񳁿��w����*~W��(�ނ����S&�6�b�?�>�( ��<k,,�P�Kr	�6�r�*/I%�|h@��*<�N�Y4�8)u�M��1��M)\+�%��_�J������@�o	�}P͕��Z��1!�MX���?��r}֚���Ɂ�'�/y�Q�ɋ葇ӅK�c�C�4oi��#d�'�T�jŐK��ݲ�1n�I�t-�\��˂��*�E��mo�zO�[��?)��CO'qw��;�_�� �y��6���m�6�v���KdEʢ=��al����w��%ݓ� R���,.�
K���'e����w�%�{˟N<�B�?�?���rD$�Z6`���`i�    IDAT\j�'���@J������@ܢC��1��P.j{�ߩ ���s�1��d\1 ��y�.��<���������ɤx��D9�j�He��.R�ʣ���Ӥ��Naw��z"�-j���w�9��������:X�8�^X�p��9V/	�@��ķ�M��|�K/1���;����{��M/��\�2>�_U��L����](	��9�\h���� ���-rÒ�(K=d ���v��W^wwy�=ɔ���{s����3�.�e���R��t% ����yE:F$��y���/���x��������Yg���/�˳�7z�@^:�2���q�SEn�<�WM�,�'�|�ƕtɹ
����E�6��M�8hGɂ����ރ�Ҹ�]�]�y:�2��E�a���)Si�5��
�_@Z՗�'mjDux�(�Bȱ�iŠ�Mq��բ@-�y^ �9�?�n @W]lF5�S/��x�0��òǺc,�r+���/@�kh� �����k��w�A�(z������]EQ��/pI�d�駯yU]�LGb.s�*	? �,B㩫+S��52R
�x�z�W��ǖ&t[0p=�} i��B�P(�G� �T�r����}������9�w�F��Y�ъ�zRT�5j�o�(V�+<���0��������ŗ�?iꔇb����S�?̓��`�=A���b8u�+��T� -B(���-��O��=��-<?����<��s����K��d�;�?@��/}Ɏ�!��q�3�=\P��ML�7���;�$�K��d{�m�l3CRV?���~�^
@�� ��?�{���ώ�K�S�bs.P�okB�/T~r�F��5u���]d/�~��;�3�?��24ħ�� �mj��R.R&:�:�X{C�=�<��C:]L��n :��>�߿�GO=�D�w�<e��i�5�!��)��V:�
P#����\RH���XHV���Xx+V�H��U.����	����`s2ר���sp�ƹV�I�5���a�A?���h�"[�K��P��#&o;�KV��)���y��S#�<��؊����c�  (�����l�[)��v�gw����u+b}�I����#�ܐMƩy��� pU��|'ʜ@$4�:X� ��c� �(2��3BYI�!P=('��w����'�H�v,͚�{f���O8�������ŏ_?��S���5�Â��v-��@3�� K)�XH_��K��B��*vt�M��f`#�7���j�q�]�p �i)�����e~^�� Y]�8��a�Gi�P3:>�s��w[AwG��T�BQ���Z���P�� �m%�_�M���m1^x�U��T��ۄK�/V�w���a�J�����j�u��\�C����:~�Oz����O�|�^ �뮻μ����j��?��F���;ڲ��i�9�5�a�o�
���{�N�U����S���"�V9D�v���1"`|]��;����g^�0����|�]����O�')�vO��Y���*�d#�	A�{6  Ϧ@�-�ʝW{�̞��VIc.h"��s�Il:�uF0o���ҍ�Ld|6^p�9���`vu���#��5bx'��k�eA��I!�݄�/��T��\p�����r� P���S
�>�\|�V�*O9h� ����i���h g.�I�k�	�gm����?�Mx�4�|��Nu�d�-|��U�(/Q�Ɍb���.����j�����l=����x�s��a>�У�)B�r[cc�=�~XX�x(����mm����aWf�,���7��T<�VV�{������8�b���ӛU�� ���X��lB62uӗꇱ1F�1��6�!���(*p��#�1�?���R��ݼ��<��)N�˟��g�.���,D�e<sQ�r��$)�C�s���{�N�H .OS�G� �oϝG�U���2��N[)-Q4���߅|�{d\j�#ߜ ����I���]9�U.�x�u���u���o\��-���L�n��ƫ�T�OgJD�v#!�X�X�:��M�S>����tK7��0!��'���@�?�B}�y��C۸��5�Rg�jL��;����+} �j����Ac�Z�j�Z�|k8���-�K��6P1�?����0?�?��%�-M����8�Y2&o��e��d��1l|��	��t�WkKO(*�m�>�g�)��ؖ�Ke~rO�_^��+Y��TRyԒa�0�H���>���[����4�/N�k��������oO���'�3m~��!�m����K��4�":(�'V��$]�]s�VѲ�]�K�#��Apw�M��`���i� ��z��d��]#���Wq�֦n��.�W'11�dz�y��f,�yF2MHC$3��J|�Q�TO8��LJ�J�eZ�C�馛�x�����9Y��b1�7�с�2����x~h}WZv�er�g�X�(`e6�5�<gbܬ��;���^����w���a��3>,h�V�#{���O�~���z477x�7�y�O��7��Ͽ���^_������W���Now�Vs���Pv9V�<��5�  ��'A`0��O�P��݁��YY��=�!��( �� :�Qx(�8������K'�i��o(�e��pjn~
��W�=�%����g��y���`���yꮲ�>��������ᕒ�C\�s�Y���1�8Lf�ܹ�������J����&g��w�1�ͳ�<�[�w�ڢ��|�G|������l����=��]s�����ٰ�e���8d�����)k$},A>� �H��f\46Sa�t��`�ɂE�͘1���~hSr�� ]�E�qh�[Z2�0�^,h�rt=�B �����O�Q����k��?���y�I�ĲG��ƿ�� �W���Jnh��}d��k�i�X�6��mW�|D%�g�d˟uW�+��θ
����e7Ͻi�	�����9��˗G������۾� ��"���D覻;�+�(>�wQ�*+Y@'�7����lyv���H�� �A"*�`����)� ���;��������aEqo
��P��>H�$�"CF']1&�
�����߰�I���u�.�ÒgO�g.)�c�PH�A� J���w������$���o[o�އ�=�3c`Ȏ��x����.Yzaw���3��(��O�x����Y��P�]*�W��-vw�����С�d`(8���Im(�_�)$��͟6	��un��RN����c����= +�-���q= �L��Y�����KA�����Һ@ֿ{���f���8ԅ�o>�Y�FoZy�V�?��5'�S�H����'D�
�WZ�^$��?xg0g�l��T�2��ֶ�	��y��=[���5׌[��s�Ps�ҽ2b�Ӽk����_i�n_ײW���b�\|�S�gf]�gm<�,�Ϳ��J������a�Pm�p�B[��D�?ܿ2F\�E�|ƯϺq(� �5k�=xE�\�	TP,��]/��C� ߮'�{*� F��d�`TA��8���6̤%sp
��<M� 
��ۓ�}���7��Omʭd��.���rS�Y����7/�q�)�?㌕E�<��c�}��~S�J@���}������XG��4Qt�jS��|�3��<7cb������%�����8M�Hl,��*�����Z��w?�Z�����d4�����¤/�I��yEQ��"Њ�̳g�>n�:�Qv��?�?@��!������Vz+nB�k����ϧ� 뎼�P9���s�I���7��������@��ͦ�~e2�s��o�{�-�A�����ڴ����sX��R?p�z0ϻ����`��"q`!���Q
�R�5�LlO���SdD�/Y�
�a	`j��P�?�x�Ny������#e��w�ːB�'=� N]�tU~RYK���eZ�x����?�wPH�h���T�>�ޟ������/c�R�������<��axfd<�_�}��˵����q��յ�k��o�qyу]]ݨy��-����6 �pQa��%`^�޽�孱���&��f���t?F!�k�Me͕5!J�9���LOr������ٹs*��wS%L(�2Zb�����9p�pǀ����Q$V>Y.��
��J �'#��cUc�B��=�>3�a�ųJy���ݺ㡭6�N��3�����g�bW�G0n(�y�7Y���(�"�L�//]�9�O������~H��+
�2x�Iz~�p(l�xZV����]�.�P�����z����s���:l��t��m�1�c}Y+�*�tXŠhT�{dUQ�-���lsR����~�UH�b�T�j�\�ϧ�rʧE�L��i��[�z���x|�N��F�
���%m.ޚ�G>7�c[��[����'�! �r����>N�K�\��75nN��"�)�&�w7�����E_��<U�r����`�*A�� ����'U�X�|�@������J�T1���Bʏ;ܟ�S��HhO���<�h�J_Ei��g�� �')�/���y�駶i얹�p�s�J����!�#wj�)t7��w����m�������-P�ޙ����
��a_�l��+��<3
�y�M���O���ȅ��HH(�\tw/��XEvvvn3f��{��/Z��*ڇ�_�`�~,�;O?Myy�; ��E�v �F�:�r�7�Y��>xܸq铓�LP�tEU��˃E(�Q��m�UQ����L�|��L�cu,_�Zuڤrְq�f���yq���.��Kyq/�	J�MN����g�B�j�\/���t��m�V�*\h�p-v<z�C��l�%p銟0^�}��Ȋ<��s��3�ِE��SOn���sJ�?��/�0�̧*�W�[�gf�Y�&��-CF5̽���ho�b�ʬ� ����q �]�_�N�S+y��DQzmy?��dXN���k�O���O<����\~��ǿ��˿�ӧ�H{�meEZ�܉��s7C!�����r]^�,0�!��e�a�;6����Ea��Wm~��_Z^V�"�Ue~[]������TAO�M�>��yYm���㓲�d]���D҂?�̼(��!&`ѽ�,�^�	�wQI���O��z�(p͸�QQ�'��L)@�O�QAA�>���m�E�06�g���4ߋB�Y�lN�G�b�#c(��z����`�R�G"w�� \zO�\4�s_��%���}�q M���p����_��| �����U�<���^ߵG��Rm���rV�?��y���)h�����'�|mCC�%����9�J�]��K�4��D�ȍg��:�hk7��~�3fL�e�F�eVL������}��g-��� ��<w�)�9(gS��~7��sdZ��m9� ~�6(�Ϻs$��C�v@�����/����(%'�r�H
Yi�Fۙ�5'|ʊ�'2�zi���~P|tO�z�q+;H�,E!X�����/�} 8r�a3�%�Sͭ�S���_~W�T��p�G4��h+���kC���[�-m��ȋ�^d8�.�K+|ݏ�j��.�3k�Y}�n�<�ӯ_����_��#��ܓ�/:�gRx��!,��L&OE�宥�����=Y�\׈��e��a�6iA;��@����<����"j�,�_֢��I�ϊ?tw��y^�Τ�D{$y��M��pĔWT��]��d�+����w�G���a�1?�ݑ�v�$4�X�:V��x�_P�T�P��QO(��K�R>��9�oX�dĐ+O!�㓬��c�+ݏϋ�p��֓�c�/Y�����z��B!�G&�%=�C�א	��UUU՞�<���:
U$*�=�]�s!kY�e\娹Ҙdd�������s�(�C{j,'�A���sT4/��Mw�W �L�%��m�ng�J�gȶB����%���W]u�'N���^E	�����_?lٲe�&���P(�E�Z(�mƠ	-��|�����
�d��
���cҜp�rQv|7����wb���-mQ%����/@K��*+��s�Y�9bd,�G:;;�^�y�U�!Qc�6lذ���/ZB����,:ml�'�S�G@�^�������ŊP��6Q^����B���M�Pn4�#�5BqṸ���nZ�ƪ{�l+V�X���}�z��6TVVvvvv&����x�kkk�.qsss��7�<�����D"1�ϩ�R%N6�;ǢQXGY����E\/%�idz�?��}�dp���ʢ��mŕ	'�Tb���;]z����P�+���TC�ВiӦM?������E�L��W_}����vk8��#�b�Kg�t�����u��7+@R���h�vԑ㶩���=l e�P����Ӡi���.g�qh=C�����)P�(-��O���֯|�+����y���jmm}���	�*|r=9�f\�R:.5���)��,���<{�g]�s)և�9����Ҧ1�J�m��u��ׯ���c��3��,Y����n�<�L^TQQ1P��F@�m�P�R)))�LP����nR>�����^����I��C�6�#�S��{K���!X��V����>�Ogg��&M�����/;r��&j�̙_x��7~���|Ruuu9�� �+���L�uG&�7�u9J崓�uhS#c�y�\�6 ƺéM���V�����ZX�x�O��o��/�~�ĉ�͛�yPvwwvv� q�xpV�y�mv�����92
`� `}}��	&��\���5���/f���\�D�)���K�i��5k����WJ�QG�{b�����I�V�y���	<>eE�{��vw�()Ŷx^e7��ʮ�3%N#E�꥕����&L��ùs�Ο��H����Y�f�O�YUU%��!(�rPQ��Ke��=hs�|)v�J��pD'%���~6S���
���s�euf~�P��VvGJ�mPS�ȕ����1��a��{�wP"�x���k��/�uQ@o�fv����R�t�u�]���N8aNO���g���[n���h����d�E��Efܽ o*����\��mI5ֳ�AEe��� �:�*���������'��(9A�O*J՛H$:��˞�������:�����&��;o��§gE�E�0�:g��M 4�S���{�.gs(Sg�j�i�e���E�p�����M����8_�?���W�"�HcMM��ٳg_s��Gg��S���1���NS%(��L��<=N8�閿K��A�,׭[��c�=����|�w�q��yvuuUD��#cU��������i�lRY�/���˭�p���|�S�Ac���x�{|�ғrPFolll8p�G'k�܋/�8�>�5��;����O��������G�WS3`BWWW�F\�@�|a�I�m�P�����o.�W.�v  �O�}D�d)��H��~��UJ��Xuu����}͸q��s	��yh�%�+�1�(h+�_ ��"sn ���[���	A�$_��*풿�8��L�0�P(�p�'|����Λ7�Ɩ���*��?Q�W+N�o\HAle�Q���ԙk �2ʌ�� �έ�����O���gd�RJ!������C�wڕ�>sҨ�:�z	����n��sK�~�g�S*+*noo��!J$H��6o>��g�N����~�K�2H[�X��&+����t_��� p"[���i�a��[��kN:餜TOj\�c�<�+̯,~Q?���xBA��~o�_���;>7�@����q��{�8��C�P���:��˗W�r�-��dӧ�VTT�+�\oS
 �s��Bge	+�!��������A�G�ic�{����lR�*ڔկ،�&����k��j���5gΜ���^k�&{�=.���#V�Z������-+UQQQ#�I�-�Lv���l�&�|7�M�e�g8Qy6B��>�΂�$�������o��7��>�z���d2�`8>��� �G֒� ˾'߷'_�&��A/)�mݸq��cǎ�rG-�ǲe����_ߵ���*p��.�+��̜�H  �IDATy�C�T���>��/�V�	$v��Lr��^A�A�	��h9� ��ۦ��������:�����g!���=�͟��g���u���S�x_����D�	�BeA�Y��=����$�t56�/碌��L�l�dM�B����S>�+�r
��M&�=u�W���O��ӹظq�QMMM����k����,)
�h��+(�#�z{���9��3f�V9�1�S�zÆ�ǎ{��X�����ȧ�x<>����wSi��1�}�qf� �A�c.�WO&{-�4�S�D�o���}_�-?m�p�)2%����Æ/=dԨe�_}������%�߁�������y�o�f�ڣ=/1���r0��1������G[_���m�c������X��l-�d�+�F)���(�!zuvt�C�Y��b�!���dk�,GnL(�[�!i4e���I�?o���ow��ߞ����[��0&��x޿W��{�ҥKw(?��������YC��h�H��СC����&�Tjoo�ڰaC���2���E��]�,K�·��gw�}���9C�2g��i�������p+	�{�����[B��F��^nhhxvܸq�������˗W�����4}��}C�P�"��}�z���^YY�d!C���}��uo���߳�dS"��������(e���3{^��8����Ic�e��m7���D"������5;�Õ�}]���m��n���Vw�X���i�<�-�յ%�%�G��F�<��G���СC?�6mZS>k���R��Ʋǽ�dɒ����������6m����N$�
��D8��ɤ�,�3&	A�d�/[�掻�q�{���F��x���a��q@�1i<�Θ4.~2N���O~�߾��"a�ya/�¡d(i��ԘӲ��1&�������pg(jO$M�H���΍w�}�_�������w�jjjD�����Ӳ��pWWW����-�d�-5���ye�%�ɴ��L/0�LF��p��<����T�B!�3�L�<��o��S���z�k����9��K`�����RH3�]��u���d2�Qc�t��y�
��P�q'��L&�{�GH�1���J$�Ϝ�e4jMd��:��h[(�t����9s����px�>}jR�r�|��i��~�`���/o�{����>ӽ_����R�;]�lV�<�8�dKE}��P�}:��%�:]��ʪ_���TD������ͻ��]�0s�ѿ'.�{��k����m�lI�w��Qm���*/-��'X<��j��/�Lߗ�~N�Iw��~u����Q�G֩.�~NU�6t��Fc����q���K<"y���!��ˉ��g2ټ�OJLI[`��j���A����mP�C����X��9�?���cfAt��S�b�b��_)��%��i@k���1O=$���&,� ��~.�� PK   �eX����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   �eX��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK    eX@��)  /   images/fdf90566-ce4c-4b91-9798-b6c065370fb3.png�{eWM�5��I�� ��w�;�a��]�kpww'@���;�>0�溟?�~��յ�ԪSGj���Qj_�q�(�p�|�@@@"  �`��롭���w�t��熀����1��
W�,��sރ�ch�!��թb���A&��A怳�>���P1��c4�{?�ԗ̈́�p�i�7�o���q��'Tj��7��+ ��x�t��5��@�4ic����}���R�&�%��_�&D�]���]f3�d�Z��4�����H�Dc��K�j���]tЋ���2������o'*�k7}���������vF��*���g�u�ҴR��FR�(��y�J.���{���>u-y)��ȕ̚���7���/��L�B^��Yz�v���~rm�$�=ھx���%����$�p�(�ێ)�b�d����RW��#|t�#ge������&$5O�v}͎��l�<��էa```v:_��(�m�Xd��!�wgKG�}p�9��q��Z����*��Qp�!S��r0���t{�M�����/*��s�OV���1����3�eȃ0 C1�H�1��Z/[,V��c���~h�~��y�o���}��!V0oڦ���\�#�<��n�����E�v4̥]���<@ �!T���x�ف&dlJà�m������b���-�Ɨ��u�(#x��)���Ŗ��7|x�Z�j�S��(u�2hU����Y��W������ݦ���Ԁ@��Ga߾�X�Qm^�{0xy���pg����w�ל���/[��cu<َi+�u"��ʨ���۳��I�#�Uc�&�[������׉������ܱr����X�rAĈw!��/��6I�˻/Ty�O�R�0�,�8*ɽM*�}�վ���?�kV4ʷ�%�Û��1��[��/uzM�g�P��_a�'y�|�1���!�cQ/ے��恑�x���w��0y���#j^�gX��n�DT}ҨL�@�"9�=H�y_`�~/*�W%�L�kH�3DB�5,�W�@?{���<��������ѻ��껀��	��/b[;��W.�܍d~UI�o�/����R��6�P�wWа,����T�^Nw�A�֪�����%����t��'7��Iy�-�r�|��cC>�܁�������k�8TZh%嘙�k�,lV3�U��{��T��}@���旜�4ӏo��g�.��Bv���sfK=s��:����ʷ���L�1����]�j���1� ��6��uj�[~|�eĔE ���^���/�O~�бd��v�z�7s�2��L��xm�$dr~�t��������L��E4O���q�~�k�9�C$�@«��
0*�9�A-p����"���A�ݻ�ޜ��۟�6�[t�s~U��q��x���}Xń��y��m2ß���É���R����[�gb$Q3�AȆb���$l��TDl��4�m���NIͰ$��te��S	�)��>�9�'���B�Ѐ��k���vgCFt-*�P�ط?eg�Y�ny���N~�
�57{zz=���a�	�ãNݧq:.�"G���-D���e��'7u�\aww���jk㷎wuj,8˚3�"�/?*K��:�%�����v�v2�1�bf(1?���4.�I"ɍǬ��^��k�N���ɢ������"�ථ�T01�Ѝ=�ꊟ��:&2��f~��P�O�Lq�?���N���r��`l�e��ܫI8�������)�,����_��K����>J��r�9Ih~yC���)!���5�н}������[����T�'�-�>*0��ʏwLx�� ���8?�|��PK��O)�I/W.�v�x;�0p�R�l˘�)ո|��,���/��'��:,�d��T������u�b��
��%Br���w?���iI��Q_bu���qՑ\�#���#��(a�t��qeg�� z��"H����l�D���b���.�ө�n��\{[A����a	{Iq&��K�vGm��c��q�h9���
j�h]��<)Iw��q�U����դ�倛j��^ ���������\���D���->�ao��'e�讛���K#��L�FPJ�p���/�_"K0v��5���h�	�80�kw��t�y�V�����U���O�Gl��t4�ʱp�ll?%�!7,5:���n�(�6�,:��F�~��%��OVfJ�z����I��P!�����'�A��F�3���촗��p�(�?T�E݅аA�F��snA�
�ϥ�=�̴�#�b�gV�-�g8����;��'*.U{q��  4E�~���N�I'���P�x��A`�*p���C���Kښ�'��O��A�/6���ކ�5�-'_dD�ۦF����Ά�()��]�KLjQ�E�~NMq* @��5���C][���pQO^x�/�-�&y	��� ���e�lYfʷ�iߝ~�k����}�6z�{t����͞ �N�qC��:;1���ަ0��)�U���vi��C�s���W�C��e�C�t�4��zp�X�_��W�����|�C���Y�å��h,q�W>x����q�������Q���Q%|u� �� �!lg]���i:���x��0�2�p��Trchuy����^@�xiy�+�Aa�N��7���]@4F�&�e��Wl��ȶvu��4��J<�_�a�n���^����h�3� V�ɏ�0����f�N���;��iu�K;~���j�۱�
���	�p�9�����Ew�'11���>{�� ����Xi��n�^^���H��3�@� `���п�jYY(��A�tޠ�������S/�:c��a�l�z9�51��ǡ	���.�ɘ23��K��~�h����~<۹��c`��.-0�`�2B��Ť��M MH�c��2�동k=��y��4ع޻Q�S &&�0����f�~�Dp79y���b�2��L<~�/״���Wz\y�-VSYؓ p��y�5�m��(�uq���{��1��c�ɓ��Oԝ��CK� �4�q�j���Jt�ru��e��c�^�Ӗ��󅤋)�����iP�rp��������Ѱ��K��9��L�����l�J��,����@j�z؀�8��)�����:����P�@��Y��+�;���?��1�p�F_�ϟX����s������>s!;�K�.��?&F2[�i&%�,ߧ��AE�o��U���n'8���?.pr|��~��"�9������Be��t�0��Is��^-�����V�k��]�������~�2����ԗ�\���I�p��Ʋ���0�_g���)�t����N��SR��O�A�O���� �A�酵B)o�&	\��ᖨ�q���?CK)f �����}�Tz�������-wfm�J�ʯ��&T{Y3�E�\r����8[�O�����:L\�A��.�
2���N�;&�i�Ut�����s�e���K��C�
B	W����n���~��NM%�����Δ	[��]DG(9��(Hs0|��T��a>����{L�d���H�ю+�S���ʅ�'$X���P��k�ζ�iS6�huI9g�TݓKև�=�w��$�o����''� �;̽��������q������أ��}�GnȨ�D���Eϭ�z$�mv��C�C�e��a.���}�î�d�"��_:|�y�,4gZ�L�1ɺ�z7P,�eT�_��h�Y��;u=�A4u�U��A����8agF��!�@�� ~7[��k!߷Qg����÷�Da?)�%�UZ���=2X��=o�5�r�+�j3y����s�$Ʈ�}��������*9��2�p�[i����~m�(���n�g��Y��v����h�T�ɔibu�3�T=}�"�MZ�:-6m�_�>G����Ↄ1�C�����Wwt�I���i��f	F��P��8��7��!z�Q��Y䖫*K�_)��z�C�r�;j��v�-�%�%�XNi=�a�[����x��Dww�Ϛ�h����Jj���hQZ�;�|����ܭY��f�
=y�ne����ֽ���X&t������.���t�@ � ,�˂�s�}M8Y���!�� �2"��>���
]��b��@�16����iE���fO��Zz��61�Dg\F��,�N@� ��)舞J�����Mm�O}ɟ�C�`�}�!�7���5it �dC�lL�$�I�@0*`Z9��2��`�x���bM�=9��m��:��?���N�X��u����Q����;�#�ï[�~#Hqi�(�O��P�w���w�����"	���W8�@P�&�u�kg���J���;�z3����{'�&.�����zT^����l2�>M����!UG7>�o_�{��r�&w��/6Ey��~��<kB���׻�N�I�p���f
�&u������C�Ǧ�;����U�1�������iDJ$�w���v!sT;K�=Տ{r���Gj�{hN����q$���ͯ��X#)aG��Gy�^��	�4 �C�	�^�X�&1�O�֫����D)�Fg����S�L!G}���ϼ(nq9�2�tR�+��eF���#؉ey>�NR��g��?��tBy�L�}�Or�:\K��t&�,GY?M[q+1�R'S�Μ�4�G�oֶ`���3����|���d�H!E�BΛ	��.������W�ɪ���!}{q?ڃ{�fl�|�J΁���e�8�ސ��ìs}J_n��R��.���ι�7r/쮎}o���=���0��B4	�
κ��ez�Pބ�O+��MMf�һ����I��3��O6����L�?fn&�ٹ�I&�)�z����= �w;zm�)�'��'|�����\���~ݚ��������>�� �=����L�o��ę�r��{�#½�o�wm�?^���]�s-7��0�B�����$���\�D�O�c������&yG˓���43�6Fcq��dUK�:4����Z�X���(��A����wā���#H2��BLΔ� �u~� .N9w������o�^�u2i�x�5�5��w��<ay4�˳HI�/��y��X�׏�II�D,���Hė�>����S�����S�_䬺i_��'a�e׎3��f�֫G	�?Kо0l$�2�4��,���wItN��f��s]w�=ےqh����o��x�@�|Q2CX0��*o(��r_^Q��ֶ����2vf�=�6hu�B�M���U��;=���s���~	��z8�B��sJ��W��w�Db%�������{��2m�ݗK��w���R����&Q,����U�UL^|�Z�$�%���d�GҫwIC���.����~u=2jc-�e-�U"�mo���9����}?�Y5��8�K��~��b��(dk���#&؉�A2+��4�2��&�(p#�u���^b��}Vt=9�M�q;�u�����S4�9X���N�A�ӗ��(x,'�.��r�j���n�\��K�MI�T�W��2�����u��uP�l�����ّl	K���a҄X� Oc%%�Ж3���J�Sd����R��Yp0�0�tXF����0E�Z�T����� ���#-�B-F�܆�?�]�<�K����o�	�$-3</M�_�N�f̊��~�x��)�Q�En��k���?ĥ9�ZY����x����Ìi�{��d�W2O&E��_���'*�N�
6�+<�.R���S�^�G͊o&BT�7���3K�����ݍ�o�0~�0���Vd���48B�Df8����ƾ��Ѻ�ʑ|r~'�"Bm����wK�lN��b�-�37��:�������h:`h�t�2}���;��-�)
6}h5���LY�� ̓^Mj{����6}�:韬�sX��е���'�W�P�g
�l��LI��g"�P<A�9�a#�w�S|��1�H�8@_�����fP��qQB<��6��
��T��I�as��!S�����S#l��}�t������P�a�蔏���un�(-@��{XV�J�@="��u9�f��6]�8c�π�n�1mڒ����d]�^�h��c�M�֤�8�f y��} ��Q	���x�^�;۸���L��ܢ��:f�$/�駭��B��,��/!��g�cۓ7���:	�%~ �J�O?��������X�sG�</W��Š���f"�
�u�t�fC�s�������4�;tڇ	�c���;B�dF��3F��
s�U���o�KE}�|�	=��9�&�Hs��|�C)���	c��*�n^� �S�y6A��/$=�N�1&K��i0�h����ߩQ��L�\�%ޑ�I�u+'���U�U���/�A/3� :Z�AY#C�{��:M%�5�-�2���h`���B���fϩ,�f�K�� Dc���	W�@'B$7i���#�yDh��IoFb�&��_B�����4�� �#�\c�aA.�%��ھn޷��UjU	,C��^��=��EU�($bP��rq�℈�?���BT�Mm�)�Gj�d��z�㦨�OzG��|��U�}�т� �.����������wb���ٙC,ddD$�hQ���q#�� :�9�1=#�Ȑ�X��Ǵűo����B����v�X����S%S��!�g�VrLo9��/��:}s���~�<���j��h�`D=W�g�������|~\��<va���|?�=�ď��٬<
?�vJ���M�C�
%�� �T�h���>�7~�*�į����ȵ�H($�
�Zn���E��v��g[�?Ĥ:¥L{�Af�b%*�����3T������G�i
ߘ�jih���&��xY�O��fB�,	n*�×}��?��V��NeV̛ X�)�S�';*:�2<8B���:&5��їf+�N����=�V���2��/�)~Չo�u�&��N���v�y*�'����&����޽�\}��O��3�ןf]@��o�VA@�<P��]�:P��1W=���k
9�����5�o���~���b��J������qpW^�W����q3D��GX�a
���9����������d�o�S-|�>KU�@/�J�t���������x��
����shu��}�h���_�����|fv��o�M���I�>SD�K��/]�P|w��=�	7U�2��mv���٢�I�D~���z}��	����g̻�a�&zF�#u�F:��Ʀ�<CHJ�����m�{�|Э��Y�f10z��W+��C�]�Qz@R'a��]/	Q�O�����Gv�k�L~�x�Jn��ʻ�[��y���bI��H�lۗ�8)ώFnE�P�U�[cW��q�y�t��S��9�"�
|X��:[��J�������O�4���d�m�7�q\K�,"y�=�T��	C��'��c�J��ʕ$�&���į��#����1#X����p�E�.Mw].�K����1���	@���87�N�'Lw!6�ۀ�5���=�?D	��F�~�	ن�y���<9f[T�	1+�b+8�m�R�JO��Ũµ��Bgw��?�F*�.\��$�x_#���7��;Yn3�j'�����=]&϶��D��ID�x��>k�7�_c |af*PF!@7S�� @��o��]}i��f?�"x4�IwA7�{y���nwȆ�4�> �.Io�&�p���kަӢ�֌2VبXݘM����X qJ������Z��=1���q/g*0{YY����;��d<�/�����_R���*�[��Vݤ�*�ڜ�fS��O�ʲ1�)N�CɎ�'�������5�bc�s��ID�Ή	�N�u�\����7S�kM�"&\��2ԥ�^:�s��b�#�po"�V'-#������Xkz��^>������FR��Ν&��v� Ix7���^�Cf�� �H����|{�	�Ce2&�?��׵��l9�^"~��o7���C���/K��~O�w�&G/��qvm��(�&uv����7{��Y|3n<�#�Ɂ�Kl������v�X���(��{��!0�2qƪ��\�C��D	f�n��_4����Gx���^&���|"�V�-�N�����/1v}ŕ�����oӉk�]Z�4����_��t�}J&��MP�G�h�	�+��4O����Zy��m����[�^�RXi7kz9��\$v��V-�>�_������Λhp(��:;�{9q]sl��wy���x�	q}���EGA��+Sͫ͒D����A�Y��oG��G5T��E�]-��D�ep/CX�H�QY6��0�ة��hK$���J��N�Ã�C��k7���ON@���,2����l�r�����p-�'J�\���9�����a��e.
B5I���â�s����.*����=�K�?��4�f;�:�׀��B��B�aJ����1V�O�)��/�E��Fmcڟ��}��_��t�l�2��.����1��g������6R�������lN2,8�
�]�S�����S�}U�@X��Ɔ�Mve;��a�0
$��P)}��7#.�T��G\��lp]	>����%t.����V���΍%+[J� �D��h�li��z�X�� nw?�x@%�>JY�x��h�VP��l�Sw~Eji��u����|�M�6���j�^�n�JH�ؿ��dbMߋ�̬�����F��U�!�k\��O	˴�͌7T����r&�m10ͬ�:�j�����ז3fU��Ѳ��W����������E HRBt�U�(�}f!�JBN�,km΂L���HVӦxG 8t���h:�A� /ɒODO;���;�zo�;".�G�,W����%�D:�C1C�5Ŀ@������z)�Ɍ�#�2���OR*dҞ:����ıd�b����t�q���c�׏��q�s�{��RQ��+�ж�mi��s	�l!���UͿ�!�
���)�;�;��Y
c�)�PCp��N�G�_�E;Wh�̲e��	���̲f���56�eV%���e1�~숆�գ��[�+�������R��h��R'��F&��	�@��8�P�'H��E��KX��G"rr�[ZHK�G)�c6R2���=n:�HU�@6��{Q�f�aAb���<��װY�O�}Q6�w*���3��#�����I?I�f��>�%&>4��y� ���VrCｰZe�|x���'Wj��i�o8��e���V��2h}���=�)O�Qe�F2�!�45�L�4ՖuVj�a쫓ρ��j�+$���L�����BU�{�^���T�� :��vYI���
-str�gv�B{t,����kk3�hƃ/�I�'�_%߿��j�v�M 3�ѓOM��D�%�͸N�������z�MD��+���z�@�wL�5t2��_~�c�E�7��G>�w'*3\5�kImt��m���~Oq(^�˘��W¤�z��%7���C;�j����p���v��^N7	a�cz��u�o�j���'a�$��%�7����fQE	6c�c��|Π��|��&� LD\������Pu53asE���z�[_�&�W�@i��D�%���Q��kA�_�4m\��T E��3:���ÄGZ	�@E�YdF���-��>?s�Iz��b��m8�#C[�-�{�뢢!t��!���R����g�1�z��E\���Qly��1sF�;/
l2��g�(e����2`�����H�Bl/!� ��ޏ��ǘ����M�c,W�|��8d0+vP�]$B�v"��GO�����+E�a&$���ћ�P:�>K�P2kŖj��0ߘi������L��o��4�Y{y^t�<6:�V��\�{�}9I~@`��;5�W���o���j�9�ѩ�Q��t���]���k��ΐ�M�7�D�_8�<�C%�[<2��� q�J��ڂ'�B&܅1{�h�����pg�-�^�Z�����*bA�ʭ
#>���+��Bn��d�bksx��x�#}\֜q����|m~�:��'U���A�V-���8=�P*���]	��Є{��9p��Ɵ\�m�ی����o����|{x�[�h����k:�h�f6�>߂����j����<�'�(k�p4��V�I+�$���L��K�5ʿ	��J��l4���t:e��<�9�PU6D\�j��m?[nNp��)�7��.��쑙Q ��uA0��H�Lm��P�ݰ`�1�ixʧS���\a�Y� �~����i����.������|�ɜ��V� �tJvLv=rq�EZ�0+�R�b�nE�G��S+o�V��)-��жx'W~�>3�_[�x�����}�}�z~�ʃ�cQ�C¤��-	 �"$��"��5h���K����g�k�e�$Cjk*�XE}�>�~����וVBVk��'UR>�S����r6����8u3�p���FM}�ԟd���d�n�m?vR�ܼ;�?�~!�l�9�������Ti$�	�vp�}�����>�CөP`�^��,��]�&=5h~�O�{G�O����[�$�G�r������:7Rv�����IF^���9%�L�;���l���&�z�0,�Y��-S:�$���f�	9�)X����8_������O����9�O�k�塩\S�m���B�+X�9�ylI0k�����C�1{�^�� ���-4�8[��8�5N���I^J6sA����ʦ����j�QY������硖�k���M�(���_/uu$#]@�>�$�!�!����Ea��=����fw�>H3�94�Q�]!g3v6*݊4������ǥ)����t��T�_�P���6��~�a.���7",�U�K:�|/���βڶ��]�y�}*�?P��*�~_1�y�.�<���%�L=�-���X���>Ҷ��*M=9��P��od����ck%��x}�ȒMP�I�]	��1mS5�Ҧڝ5O�`L�@卬F�
�%�����7+Pۣk��I��,�G{4BI�0�1�֍�.�K��~��h0�4�E���;˺�~�{����,S�Ѵ��i��=���.%��o�˹�A 6��Z펩��Í�ݿ[�q���9�$M��<q侺ň�����+���������=ʐz~Ffu�X�|�?��}o��K�!p0���ur���8�lD��g�T�>�P7�����a�"3d�3{�
g�������J��%�����|�_#��N������f�j�TO��9=+qT�6�#�L��vf?Rk��|��g���qm������O{�֦<���K�ڝ�E������(u��տd�!�ӗ�A�vi�d݇����f���i7��тG��C���eCX0�h݀��A����'^X����'\�eP+�θz��J��A7�K� u����S~�Z4)��p�W6 �����$�+p�c����`&X��8Q�p��w����Ϸ䠊9�6���A�H�ӗ�u�pV���*}���F���x'�ssd�����1c���{�L�z��R"��o?E}pA����򩓲��Cʜ7���*G_���cv��U%[:٣����|��&��y�|����C�w��fv~]��__�F7H0���$��p<^$��E[BM8�NEG^&�ht.�C$�Q���l�uo�޺��`�4iM�w�q�j���cN9w�5u<ǹd'Y:��n�����.�m~�}S�֥���������x5S�-K��y�����5]G�_�R�-��x`P�8�v�(O�>�n�ݣ,T�XQ����w��������� yR"Y�#l5��`_��ݍغ�G!��f߅�jV��+�����ƴЅ�����
����=��޸ �*
Rj:m�z��>�XS���=:��uy��}F (@�ɽ �X}���p�&Ϩ-��a~'��J�'�:�\}NP�U�&ֽ�m6�n9B�����Z��+�V�[�=���:&���H����ʄ����wR--VX'����kT�g/S��*9 ��T�x�r�L�����J����#v�j15l��H��`����07��gQ-!���@}U��#ƽdL�6Ά��
Ȇ5��?�k�2C�r\`q՗]��b�w���t���yb�h�&`�!�+��k0x�í�ϛ���J�{[K�x�(u�J�Q���j�8q��j��@]"���z�8e�i!�#�Y�Y�1[C�u(��| WuFR��}�S�-�ƹ�0���Q���.�6wm[w$��Z��C7FMЙ���o���ZTnSfv�-a��i\7�φ��_�v��i�u,�eV�;�'ᶔ��B�	��s�a��5g����'|����%���2��\1v�Xk��_G��!��a��H�`����*�41`�~�u���cɈ��t<�	�b����a���0�$��e'1ί���e��c���
���fjg�*�c-z���m���ٚ�����a�fV��ߏ埞�7��-�cfN ���ˊ
��C�+��a��Ѧ��#���a:=i���ݦ]�W�ú�{K6����*�%��d���.�7�y3����-�ʸ����G*��N�Ѳ^�����}L�[��
H�9e���"#Z<��
�F9�6�T�B�ix��P�_�3�̪���W�f1[(��O�|�S����|=�$���b��X��٠�f���:{��J�p��j~��,��-ST�z
=C���+��}�?����X��-�H�k�~�}��XD:I��
�q�h��Dj9�+#D��Z83��På��{��K�?@݂�uq���Tȟ<���J9�!l��|�3#́T�T N_����"�4?���i������0���`����1�n�=�����r�(j�!H^�wp�e�<���\����haBxPXFiY%�Sgd�����f�*�ZH��ɩ2����tƩ�*�(RU+q�h��z��h��/�)ݳ�P�c�SPs�H6���i31�~42�x�Of��l\,���\���x}Y��>9=q�ґS��U�.����<jK�l���l1�#�������m̲�����X��u��Ē�)'�Y��G��}�e�����ū�b�3���n��o�\�G�wį�/m^��P0n�ө\��r�(/~�=4,��.�姚�LCn7AHB�٫~�#�y��cl�qt�*����ApCZS��.fe�s�6������{��BO�<ae:6텖S��:��N��.�Z:0�ͣ������o�(O�����'��f�y"��8���M��q�U�<X�^���>�!R��q��<������z�V�2"���s0�_�5E�HJ��ʿ���P�,5O�!��1��X��7Fq��̔$��j3��w� ���k��[
7��<�E�Ӣ��~��x�B
j�y�I�.yIl��}�-ɌNR�?�$�
�����&LC�DfP��R��J���݆�׈O���Ά��/���,[k�R�yEaQ����3[Ҕ�ڪ�B�l%n�k���@�K��fT�
��ٗ5G,H�ߴ�6r4�id�LB�O�[�j.��e>��f{ġ���@�Ñ$����'���䱳�yl�sZY5��s���5����k���7{� �c�Dqn�C'�q���Љ��S+)1�I&�4W����+u�8D���w�ʴ�s4�Dse���;tQω�{!H��$�����n��P\��n�y�m?���Z.�
5���%���+������/�"Q����K�K';�0+�O_���fpm�ֶ蚾C[%X�Fǳ�	��k��p��/ 5���Ge�K�;\�R�+��2)Ʌb�S��&�kS��R��%>Y�'�M������"��gֲ�����j,���<�K�p���Lz?���(�h���p��X���[zeON��B���J���qSZ%�;/SSr�A��RO�>�g%*V�9K!�����,�M���F�� �ね���ѱ০8��r��wa��'g'���km����G\�Z�Y3:��#�Mp��I��)V�f�֨���ˏ6�z�<#Y+�3�=Z U��Wں��-2⺃��>Ur��|֩^n��n'�Io��D%	Nvr���f2᪣�L�!JÞ���7����[����̖�����SL��tGy��i~�Et��TB6��O�Bz�-V*�A��o�Nb#W��J�,�W;�EZ�h�~-��:��
�H9��i|�
��󝾶Lw(a�x��ZG�(.��<� _�;dּ�5<�?C6���[�D~p��ep"P���4\a<�|�E4��CLT�Gz���P����6~)5�^R��4+�{Oc�m!��U@��s��~#���Ygw�Q:{ԄDA�Hǔj��`�l���m�z�T���^������(��y��yo9(^<iJؠ�X�D�H��~3{�Ze�hz�A/��ܬ&�L� �q�} �#j���U�ea����m�~c��J���l�
�R��3U{��a@ej������7��U����~kz�j���vi��&�h胃F��%=��o�ETYB��&F��l.<?�-I3�t�'aV�D�^�$�~ř����闧U�p�$�d}!q>ah�Ă��~t0�jn����#��)��Uqs���B�����	RH�	Z [��������U�;Lq�t#�*��9�#gCp�mX�B��bj�U4��ݏgY��,�}PZ+���OZ�YMh�l�dH���c1�]�tP-����
�jQ JAq8��|��Ҡzc�Gh#��p|����2�b���QI��H���;
W����	[�e���ALK-є��|�L8Aqrp��s岎z�B��5�Q��0�b·��5�X�H��w�~f� �i�p�Y�~�.ஊEH�4�/}�J�hu�[��1��k/o��|�ߊ�d�cf�AcpWq�M��oJJH���t~u(]�ݚ��F:VV����GL����4��f��'�������G(=Wa��?��)7���`{��P��s5b@ɠ�4	�03��+�߁�pߔWH��^�M%A$^9�>�L�o�NEt8A+�=�?1M�}a���V����ϥ���l�'@a�dI#����h!�H?�M�i��Y��Q�m�y��Sx�%պߙ�!�G��0m���ɓ(�B�n:#	ڹG��$γ q+�x�Ɋ[dO
�)�@y�>yS�-8.:�=�W4�k>�f&NWtO`�^�57H6f25E���vi��4���W��Th��� ���eۣ�ub��h��U�7V�7j��kc�{u��M^Ou����p��}�S�t��KSf�`+�5K�F0��G�-��ݴ%q����2�P��I�D�����-��?�i�j��"�lqln/aQr��[���]�d�XL�B�O�H�F��ڽ�ϣI~�<�H�8�q�9w����-pcRފo�5W�����6����y�_������yhiu/�pS�(WQ!�O��hn�@���r�|�U�Vfٛ��!�㵪�R�+_���6E�f"8�i�)bR�w�p��X�rҹ4�؋�t�vDU}����ΆCo��#���X:#9�.�%��7!��W�d�q�Y�5v[&!�/6�a���&�}Me���5��\�a�$�K3�=�Z��K�y|	�x)v��3h
I�k�8[���CY�9�"-��b��ʲ�8�!�[�ed�Ρ?[��m�gAX��Q_2!�2]+�*�^���_61��ΐ����F���c]׽�J0��;ad��n��|43X�����?g�/r��h�?I�tf���X�f��N7�i���:4�շ���T9�Tɝ�l	�%��5�J�@ա2Yg�t�<ԕL��KO��W��|І"Q��[97�b�;V��K��F�]���}9~��-�
E�AЅ8���e`���5�K�5T�-�J
�� ]��wE���d'�X��Y�{L�Ͻ�/��pd��Х7��ofM�$��n7�n��ƒ�P���z���6kjMx�>!�O��G����D�����do�� �����}v�zﺩᩋ	���=�05s�T8��x���T%`������f�P�F���1���i%�˥�9�`\�&�����Y�s����S�l���k�t�����|rZ����$7���"���C ��	�]ωs+5Nf����0�?t�k:�V�@j5��泥������hƄ��m�"ywc������N+�wa�,��6�9c�%��J�Q ��qx�e	�;x5��������HB�	���$��#*����v�յ�?9"M(��DV~��Z������N�^|�k�S�B���Ch�0�'�	����ŕn�dc|��`@����=���p�NkWm���F+ox�l���@����U=�}�Q�7�I<�`2��� ΑI�R�e���L�J���gA�^��-�ˆ4n��O)@Y.���߹�*���?nnl.���,?w{�e9xn�c�#�g2!�����ԇ�p����� ���֊g�n6jg�ݤ�D��w�k����<B�n�w��ۣb�=��K����O^X���+�.�L͗SOYf�j) �"(�����3��_����L>t��aݭ@����_��X��?�Vv��Y� �\r�B=��u��7+_a�\6�Z����oy�{߫��I�r�����{�<��	A^h�ha��,9Nλ�U��̳����m��fx�^].�`kq�{��y�{6��	���4�!��`��nيSe剧� ����|ꩧ�� ��yh����Zy��U�c2���7�?�,Y�D�z��������؈�E���}W�k��rQ�Ni�\���0����faiٿ�[3xӞm<W����v�1Md�̦$b��6Ԧ @������ܢ{d��sn��`�{3���fdS���s�|<�	�,���eB���mA�&)�x.6*aͨh�����Z���7�n	c
@םq��N*��e��?��I������#��r���m��B%��B���=�a^LJ�l �!����ݽ]
���B\�L�=���fM��j�a�[&˫/�B^{����PA��)�����G��C�ۨO��c��>�6���+L�I'��e���Ym���������a޹���y�0  pL&�(�ʠ0���c��]��ʕ��l�/Z�$�d���+�/��dD.�u{�r��%=��q�O��g�cNF���C悈�2��m���0.S�k�<��s+M�j���)`�`�N2V�"�9Y�Ƶ&Ș]0�7������6�8�E�(x�
�;��m��� �� �XS������/lIg��m���e}gW�(J-f�H�`�H�b��@�iZZ͝�/�5����>�Y�H�U�fLozӛ�G?����|\(8�:H��A�� 
a�1΁�q����{�9���uP�9|ͱ�&n3�!���VѶp,�t��Y|��CK�a����I���h#�YP+�y�+����ʍ���ovъ7�&Յp�={�Q�^�8�S
}�R�`q[�V[�y� �nb�?@��o���<�DW�[锉u��D+�� �mj�Ԩ)Ad�\ 2K�K!�j�Ԩ�ٓ�������S��B���jx>�R�pKoP����s][n����砐!S���r��D%��Z&ǘc;�)hf'�E%�S�;+0"���9���)Ӎ��Sk9�N)�ӎ[_c>3 �$��U�Vi�}��>4z0v|��|@���AK��xZ�ZV¬'Xp��M$��Z����Wf�c�!4�
���`�3�`��orB���I� C kD��=��D�Z]0�0AH�:��4%E��9��&S���q�>���Ae��4Z�ʲ����{��[�Fv��l62�X�ڪڭ��S��؅3�5�	�^1�`Xd�7k��[���1���9q���q�ݾ
��ϸ �}n�}U�c���?X}�|l`ι+�"�u�jSxP萑��\�����cxM*9n\�֔ƋB�D���*�V�}�>G���(u��.>$UyAY3߳f��x�L��@�(iM�V�y��k���Jv��M��.�}�z�ɚ�w/��:a�����^˶`�c}2>B%�c��H�A�������<hR�YK���Cca�F���# Ԣ�_e ��&:M^jVdH�	]F�����'�9�	�&7L=������L�Z�ٔ�4�8���2y��j,�}{wjuC<������c�\Ư��76��zfI�C�ɝ��(�x97�;6���q��Ժ����2p������$L�q��]?�мO��.�A���i�3��j�T�sq� 7��bl���3�q�C����z�TɨR0x��n@V�&ok����3g��!FѪX�3\: d�gRz���ף��F�fQ	����Ý��|Í�p쨔a����G`n�t���o� �7T.�4ak���ΑF��e5@�'��H0X,$�KޠT.EL<ה�����ӛYtA�ܰ*� � ��P�Z�|h2�Ajl�ri�R��Ak��1Q�@��}�?]#��
�4�kt��*8��s5�cw�i����� ������OF�Vo�68:��}��Q%V��;wFnBׂ��B�G�w�n �V�{b����.��2=� \�َ߃\��gD	�p=h�(3 !F��Z0xKbk� �lT�G�؏�DH2/�����*3�Y�ZdAֱ�����ڗ��S�k�PR%ݳRƒ���c�*@��芳�����z�5:�pc�0���G,�`����	�*�q�tsj6oh�R����M�h��z47DD��0Ml�FZ�į� D���8��R��@.�!���q=�H͎.�Lʞ��&C��v,۰)ߨ\�ճ�`��i��/2�t�X&<����oW�4炕S]�>��=�c7�t�n>7�]����;2N0�~UPD���
��Z�h�1F�}�_q����~��������8'��abS��x�-��d<\fH0��,@�0���	����������߯y�k���>C�_���� � 0@�l��Z/A��6��BU�޾^�_ 6
����V��,4�?~��(yYM��֏����
E9w��7ܠ�?ʺCQ���
~���댖�Zfx��s�X��`L`���q�����f��v����L��f
_A��R��B��G퐈�������Zh��k�>{����]��ɧVK�*}���Z�@�YlQ�ޫ�G�;�O"+-��.4-)��) Z�T@W��v�8�Mr�>��`=@��&eB	���q�\��K�.�x7(��+�g���!M����`�{隵�ۼy�BfP���KK��up,�{�'��\ (`�x�5e�b��!��KZT�:��"����F��{����u��S�į�_��g�2�W���rkn�"�g̷E���ݣgq������ *JVٲ�����B�yC)g�E8�T�xp��+�d�a׭��v��B��1*M �����#�礹Z�;q 2w�(�M��Z��+�B�ߥ~!��ν��COjUO�=��%��G�n]���f�$5Ϗ�:�7k�'�#�%������_Z�{��H����6͋[eQk����܋-��$޿�����w߭��:9������&����`ʌS0���Ƞ/��zX8�t� ��f�ƅ@n^������,�×���~���Gq,�����gsv��p<~ñ� �|�I٢�O3v��B��(@�U�u��SOJ�-Z�y��ǩ+4O�e�&��0 o�O����[��`�"7�H�����q�� ���`��S
�M�Av5|��r%u܅� #�@�Ƥ�ZRm��=��<���mL�Nm6�|����n��֐�^2�-���������� ���F�]�IYa��H.0B��B7m,%-�e6=��BW@b79j-6�4��z}�[%�;4�@�k~������� � ���C�	\�0?���� ���r���eP��Q?� 7�k�cG��!�tAo��袱L�U��k|�\U$��2o�+�j�{�N�/�F���	_���%t�Kk	h�����0��ZP�h�q�k�`b"������Bak��?��gRҹq!3�B���es��@n"�L��Ԉ�v�b��ohz����ק@�����\��B���6��w�N��]Q]=V`�B�n����_ށcC��9� ���h���
 �#H���g~�_����0��`&8�����Dt��."ąC2�ߏ�i�L}7�׍Q�� ��pqshE0Ǆ�D�ؖ��h}�0O�/QP�s��5�ǔn�1�u(��^`��5Np�:N��3Q �|}�b�� ǂ�(c@&<��ts<��606��/Aᅟ���TF9wno�C�	����΀�3qӻAN,.|�=>mdsp��:l���.�:V����W얖f�,GG��� �y
}eim�&۷�UV�Ug��:�4�7�X&b�� �(�_{0&OA@���,��l���Q�%��5]j�86;|��3�b��,>�8�b�q-�tuv�0b�<|��l:Zp���5>��I���q< ��d�8����?�=��83�)p4���\�ŭT�ZXcO������9{Y�v=���B9�bE]�%-����C�K_��&��Q����z�9@�C_|����q��P�y�_��7���+����omrq� 6}�4��F.$���k��(���M��f����Ѓ!U�[�R�5&j�4�=X2]ʅ�m�e���Z�X��*�Mii$��w!c���3�ʶ�.���w�[�����I.y�7F�}��`�6���\p��Ua�a��
��[�S&������`� O?1�y�d�T�������k}�k�q�x@�L���7D���Xo�jH� ��J�lI��1
$�V��gl �#Z�`�e,�*af}oݺMv��"�]����݃]M�R���e
J�) "���泮C?���T{���\��J�Pֿ���u��O�r����:��?����#C���T~�\<.' ���+������E�z(��ڵO�=��J��\�Y�[���
T�D�K��֠�. ]L��,uiycMsHd��w�� ���|�)2�?h���oFv	�
����;������#D�v�✘&�����*�87�F���:��lὕ����c�7�	��V!MW_}�Z@���q#c���z�*���O�T�&ċ�̃���@ny�������2�I������c��@c?[��{�V�\�x�\|�%�kj�b����Ui��|�H�P�����B?U�NGx���=��c*�+7��E�h���Z�J���*���\S-����~�'���#��-�j���6Lm�I\<�\��bc�*	Q��N^5��Æ-Is>-My�8У�/� �V�`���m���O���>�}AK��A�:܅ձ����/��PD;L���,Y�9���
,;�5`l4�/���'�|R��c�6���~����y�E�
w\��eR�V���$��K$O�m�����b��\Q��н�w�Cq�����d\L�" =�� �YXXn�9 ��3�0��k����.����|�[���Q������/̾��%G��_)�TE B�GU�T�E:���}�,Eb�=,��P{8�󬲩��la78�Y��M֢�2���������9V˼c�����C<(�^\�%f��N�+t(�2���ɠ���'/��n��C#hmn��^q��^li�k�n)4o�0P<�}�4����Ȏ۴�+�}%�fWC<��(��ۆ�]�2e_q^%b$�p���!�l�fq��$����+��@Ҿ�V�,i�(�b�����j�Ę��4��e�Wv#J�>�'Y� D_4QR`~``�`R[��8n�����׍��w6�p0OM�:��A��q5z� 6e.�U�,m����_�B	��Gg6�j6o�$�=�Z�Ο#���&2}�4Y�dQ�L?%��T��L�h j瀝~�{ߋ~�~�!��@/������#Z�T\p�w����)p\���I^6cW������^�sF;���(H���=��@Qjn�*�Y.��1�A����\�W��@AT ��c2�xr�)��+�kk�Ұ.1��vݻX3hԂns���u���e,�>���eR��C�\�Z]WPf�e3[m�\J�+��P�y�3���>ʲk�G��k��FN;����rQ��:tĚ>}�E\��`B_w�uZ��6�x �IiYpBt�d�1���k}�|��u1V�}�g2ZO�%b�� #�����;8��e��k��$�*d� l2�M��%�nj�����K�:JD��&r���w,Ǎ�!��H����(p�(�+������[*J�P��x�jts@ns<#��<�PD����V	�נ["���-�� ���};d�]j�s6�f	޳��y�	ZP�J���E(8� %��#d�z��}l)��ZO�ׁ9����#����R���׀򁜌׾�r��F��۩ �fË�v���5�'g�q��6�w���$�,��Ϳ.��g��d�Ye��^q��r���F[��"۷o���{��Ӻ�ʁv�9��Ur��ʹ|����>�#��b�]�9>Wl�!�/#ӧ��Ν�d���֔kֆ�U�Zj)ؚ'E���i2�Qb�fj�����H��"p\+����S�fi����X\+�����x��P
���j��j����V���g���XC
V5o֕"���	"���ȃ+}��``��`~Gȧk}��4�9V����B��92T�tQ�X�:��/L�4n乂����VY|�rm�R�x�W�\�I���S5��dI7K���h������_��_���B����&�ʤߞ�EZiHXl��񤣳W�|�qy�чuMa.Qtn���SVi>;���<���Rr�D�b��{�?���̀	[�p��y�*-�Ma��r�}��R� K�_�Z@�`�c`����m�������vO �#,5Lm�f=�7����yg�M2w�B�>m���K��κ��ul]r��À�ϩ�9�?�I�]�>lb�3w�2a$��Dl����1��A7���k-���R��V?��ƅ��!_C��HVz�pu\���� �u�� (�6N�r7�}���h�=��w�c=:�>6n�[9�*���g�]��D�j��=e��*֌��ڦʱ�N5V�d����J;kR�γ��E���S�yGa@X���1�p��1c��-�o�p1G�c��Ռ���J�7��=&;w�0����m�7���O?a��.9�3����SČ`Yt�t`�;���h[�dB��x�J�	�	�g�9�x꼱
:�&�+�}�fО1��+{�w�r�u��	?�St1���2W�[���Ѩ��|�fvw�����d��=�չG{���,r4}�ثha�r��c��m�c�	ƅ&:�h0����5p��D0����̰9Yր��A."��&�t3��Aӊ�@�B��tx0��	 ^�&�L
�=Ρn?Ϗ����ʡ�?�!f{��E�!KL@`�
�O�����H#h��$Jh(ˉ��D3
Z���Ǟ���}.��1��P֘@���f�L6L�j�)����K�h)���z��%��,�[�����1A�Cq<}�c�X���Y��D�pЧ7(w˾����m�Q�ɓ��W6��QZ2���+=����+.����Y�Dݍ��)�!.���'jIg뭫C�M�F�L: l�s�����)��z�̝�n&�7Z��P�����}���
�Ǥ��؄��N�5�&tr��sf1���H���0�L�f�I/V ��u� ��0=TJD�K�KA������e�����S2�K�/� ����7���������N8A��N���ʏ�# ������=�I�e�9I��C����o~3��Z|X�lr������k����w�|��%�i�����uP@Q,��}-�u���J�{�U� x=�����X�F(V+���f�K-�ַ�U_�������{J
�����Z���:�%e��������M4_~oo�TM���^������[.X,��:S�S((�z���@�Ρиg�A�HPH\�S�LW�	S)϶jKy%�:��h�6�J�5��.D�{dR�$ٵ��M���Z%69zw��t�x��~�^�E����NYֲ��im�I.m��r���E�R)!���o#��Z! �XOl6�Q�o�� >C\4�0@�.�G�+��:0Y h���+TS���������|�Ҙ6�]���2�pʤ�
�۷�h�}e�+�����w�B����5�gd)
�qpO`T \�)��������5F�s�O�	0B������
��A�J����j��]pġ���d�_��v�/�˥�2o�!�cm��P4?�s`�̜�D�F�+�i�T���s���SU�?.�7˖/���g�8m�Ƿ��-:�_��Wt�1Gl��?�vwȚ'�ŋ�Ȭ��e�_�4���^�3�=�roi��Ï<(�/]a�grdMn޼�Go�3͢��2P��ф3ƎZ��93�6��l�~�L�fi�e5��VnՒE�Ф#���7��C��\D�?�zܐk-mi���'�o�M�ךg(X �{��- �?c�\'1���h7!���nA5$>Aಅ#}���c������������$8�52W\��MX�((x#@��+��2�� 0Pi��#-���&����wn� �k��q����_/pK��ѳ�>��G�"�@�k%!��6r��D:�@J"�@a�u���%+��_���eS����e��Ge�	�$�d�~�(�j�%~�C!¼3~��}׮
���AX������K��	�פ�:��;�aƻ��ת������̄�
%��n6s>$
�:�q0~�q��=p��A�ɕ�If�E��[�[��,��#BX��Q}���m��_�����;�!g��)���m�ҴԴ�=#T����O�T4,�(�,��%}蔟Ua�����C��J��)*:�p(n������}6wN�4vb��2x���، ��]�	�bW��0��i��������<t���w��C����Ѳ�𾨀pL�}���;��#�{�6D.�����8�pq���RPQ���g�\7���<����p2T#�3�M�6���}u�jv���X�3��N�9k��q����[Rf���=���c�v��U]�{h��Gy$Z[ �0���]�7�e�+����	q,V�| N��b��?�y]������Z�{���}��0���o1������f5�b��S9�M[,9
Be��S�<����� �!͙��f�h�A�*�XHnh
�|.�Bɨܶm՘�״��V|iknU���#!�h��Y��|S����3���G�K%V�g�?d.�r|>��*�4�[4�-pr5f�,1=O&��{@.�хK�̏�w�%�(-���Hp��ܠ,����0��ɀ�c�2l�QQ�x�i�1�D.ѺaN��=����C#�K����@ �4N�ux2Z�1�^��a�a_@1*h�W6g��t^�����+�j6����X`�yͫ��y��A���,�����
���w��	�
����
�2u�qъ�eZ�Q���Y�ip9�I+��9s��!<�2�u�憛��?1��PD7 &�����6���=Ř�U��U4@5%��)��}$PuHW_��Ɛ��877]�(I�m5�!x-$
�ǲ�O|���1Y��t����b�5�͒�޽)�z�t#Д�2�`���M.�����9�x�.��ޣ�&q3MyW�e��������Em��Bf��� *�-��
>gv���;&�1a�P@���ǭ��<�D����/>���?W耈v"S#�g���
5�1�C94���*a�J���߾T��7J��Հn�Q�̝ky�����29mʲn��޿�Eo�EF!	�f�z���h�Y�e]��.C�M�k>���=�ܣ�/�ti	`<�Z'ˌYs/i��gsm��t�î����Im�F �x��3T �,��6�����z��?���v����}{�q�d�tvwȹ�](k_xFt���KS�h�d]f�m�$9jANҹ=2g^��d��ps�Իꪫ���D �����N����(&p<nb��&�M�����}��K�Lj��+����V/�@$bf����"�m�X�~4�u�nj�.4�ڸ���.��L.�P]+­�J���&�1^� �fܺ��5;W��o���� �����(���$өU7&�rqc�u9NC) |>�y\F��	��0Ǆ��Ұc^��B���R���9�|Æ��q`�с���d��^[�Y��ß� �$�L�9��0!�hˈ��4)�w�F�v�ؿ���kUY�AY�9>�' �~��� . ���K˖� [�m��[v(P��y��PpSk��O�5O����j��=,��>'�]���R��~0A�>���<����<��cr��UƼ�&}=�̝�H6o�&���/�*2�\�Yc�Z�ȢE��Y�\����{�N,��/~13�.��ԟl
bLH���vh@��~.:5+添d�ֵB�O�u�����tQ�j!�]MS���tv�� ���ʨ�[��M�'s��7�C�k���A.f�ǻ�DfF�h�E�Z_�8�v���d�|>���j����
@WP��Mܪ�'�I���q��߱E�`;�]��q�R�G�%�g�[!�E*���3{��s�z��^:s)�?��ޒ���<u�t	�e��
��ɀ��Lׅ�Ak,��)Dρ����>��ʧ>�)��~����H�s݊ p}�֚�|�lE�tv�ɶ[e���77	�VI{n4�Q���'���3t��ث(���r��R��_S�!.@�M�[o�뮽Fʥ@��Y �k!V�?��J\$U͘1K��XN9m�6�����[�zu���O�G`����Gsh	`��>�� ��!& �VS{��r�@�y���ӹ_U�\�G�v�����d�
4��2|�h�hM��ۀd0��.�k� 2
��e$W@���x\���s�)��!ƙ5\
W�P�PP��w@�_�}��u�D�w�X^�.)

�q�;D(�-�x�P�k��;}���U���:�@72�0g�8��W(<𗷷O�Y��j= �����E�Sr�+��+�`&�X3��в6Ϭ�q##w��._�ׯ�1�5�\�l߾�X�}�}��������z�{߫�$���]:�)|���_����2c�\��.Es�<����#΀�����rs_S���+*��*R�DP=���o�3���!�U=Sv�L
�&!C���.��~_xѥ�?{oe�Y��>{�]c�IwzHw愐�aPX��̹�8� 
.��\NG�\t)2xQ��W�H!!�$9@�H��t:���w՞��{����U{铳���*յ�7��3��ɮ|���A��� ��l� )����[�����1 �!���x��b��w��k<��M7ڵ�^�X �!�.��m=��-��up�+;�R8;&���%l��Ш�w�;x���-��m�52���aOeSfIZ
�Єc�^�ȩ�6ŋELD�DL�	��]�G�2AYeo��@�*u�T���!b�F���k��*Z�&5�Q(c��)s���i�e3�B*u����F��Ԥ��9�R��Ɲ2���'ռRf�k�~r-��2?�f������v�s.�|;c^Fs��9J���9i:�j��y^��C���G��7�ךA��מ�y%�s�yf���J��9��V��V�c繶�����x��h1oذ��M@�*A��_� ��mp�$�~�sx��\?�?kn\)U\�'������>�r���V�6�\u��$�YPD�	A�B���W9ae�4�O|�U��^�:_L�߳I�� K��ˎ��O�Uw�Z �� ���čMQ
l F�{[>��NMuY�)m����("�
����~"��k��Y���MoT-�)������W�kP�y�G��|�jhb\O��y��R�M~�7�c=T25Ʋod��
�@(�c(�bl<���I���¡�Oe`�!a� �&��0~1.�Ȼ� �^x��)�)�nP�}�	s���'1<1/�m�w+�5�)H4_�#�d
�;��(_�y!g��@���wx��pN�A�λ��]av�����	�2�hS��iw	x+���,�76�s�O�B��u��(M�g�p?4a!H�W\�_G��6m,۶�[�λ��3�mb���pѿ���v�|�8�,*��}���
��b��O�?����ߞv�Ev�3��o���i �$p#M�N>S�3bʂy����ӟ��8t�v���O��o��661ލ��s�p]\���z�T�{eh�U���n��׵��J��C����an1��.�A��.˒b=E�������!'B������pec���k^�':hD����P�5�%�=ER .��'�t!|��_��\�/|�δ�u�J =/{@8�t nDm8��Ĉ�׿�-�})���H��`116���B.?)�?��Ow�������b����"��\!"������'?��o}kW�L5+�M���LEH2�d^ٷ�SjӀ��¼0.��QB}���|����Ks�&��<�&�Q�{�~{��;7�fZQvdHs^g���N��K�p�g'�F)H�Յ�Y8#�S ��d����ǆ�ne��h�n �L��?�|�㡞�x�A0_���&��0¼G���ёh����u_�[o��g�$ʜt-�������������:D��<�h�>_Z������i�س�������wo���ZR�zh���V�~a�F��DȦ�T��ɒ��*t�<]h�v�i�>j{�;<;�\` ��o6�G��=�K��@t�Z��7�Ϋ^�*�w���*�A�%*VyOȑ�F�Ď�Di�H&���qe�� e��3�xS���D8D���!��nਬixaF)E�*ڗ{!���Y�� �C��<�@�#y����(�����B��W�W6\){?�a0A$<${"��#80؊~���=E�A�T?��O�{��^+^bh4�94	4��%�u����&�>�\�T��h�t\C�*����&AP&�ά�C�e>髊�@�`����s��΀�?5d����<}�ޙ[�瓋i�����?������v�3.�y��.4�hƌ���Z��f�_tG�۲�ϱw؇w�xR>��}�s͓���P�%�{�� �� ��D���N�CoP��Nx���uVe��$jB5�i^uhI�i����\��o~�C�!<"F��H�z���F�պ�a(�i���6?;e����>RN�P�s��	�-d?�������AܐH���7T#��T`	6>Ă�90�*ϒ������U$Z�	� ����1�)�"���4���B��Y9�"�����
Q�@s?��ϐ�d���B��{�~q�G?�Qυ�Drg��P�����{��!�H��)��!
��9��ClIj�X�]���ų��r�i�ar�9a�`�h*F������u��z��_�-	��2Ϭ�`42�0P�
q���_�����m�Ͽ��?��cR��kVwn"X�f��:�<�X�AVd��\J�� �V�y�~T���ce]�3�XWi�eQ�W='�j4f՛��꙱9���A��d�	O�����R��O\������K��n�9�HNJ6
B�懀�i{SW����������o8����ol
�8
�d8\��9x�"�mi�����7�CL!(%>��!=��#M�BAuVrۈ(wp/s1�:$q"D)�5�ZE�
��D��k<�k���@���* v܏���X_K���a�1	P�;c�Y8@�t�y/����ғ�E�Y5�-�*/2��nC�@�PY2�DK���Nt��%��w40�>c�Bg.y'��0�Y��~�E�+h|��4h^�	L����ݚ=�c i�B��ǟ9r��*�! a���:�C�AY�琺^�h1�s��w��?�A"~�7~�mx0`L��%�F�)�UB{\�����#f����M��'��N�6��I���I�"�r��>O��xD"/I���&U�������~[D�JQ�,�!�mE��J�ǉ|!@v�j���SL�u�!v"�����|�c�C���5%oh�$�8�X�9��Op,��1�*��sH�Ż ���x����,�i]Fb�R5�hD����^������@Ӑ�esк�/��E����|(�KP!��Ar�鏘&���i��^�W~Z�]9�i���
�VQxDI�k��\�c�b��aj�����p=�DJ��h�p%�;��jt��Ԗ��,��)���t"��V7�R��4Qf[*G!�!g�����<���c�a�s�s����5ߩ`#�I��ƽ���L����	O�����_�Q��æ����}`%?�^UL���>Tw�y��*؛^����R沴EO��/mz�p���ik�w\+��7iK����6�s!����Hlh2��2x'x4� |b��$m��8��Gʂ�+H�Z{f��:�`���,-�#y��� ��Wy�@�U�F�T9�0�a�r�4��B�=�R3�m��N0U�15*s/����+*M��҄�H�Q0ϡ��1m��	舾2F�B"%��&,�Q��#/zFz�41d���\l'$G+I]P%�����t�]�fUA`��|م1�O깕/�܈KQ�V�a�SGm<�{ͺӲ~������u�7��.ɽ���ޑ&�%��`��~�<	�Cc�ӂ>��M	�FZ�[�Q*,�?�'in������{��S�L�Üb��Z�Z�Y����\�����,I��z��m��Al�&g�!�gO��A=B�a��*C��(�=i��w|b�_ �0v�[��C��MQ��H�u!L�7��	B
T!�q��v �0R����4 ��3�:����-oY��h��5���g]B�W����p�.A��	��W�
�]�H� <����?�o��R!-b�3`���	�]f��[����L���O^6��Qqi�3��G�G�W��H?�%#��ɟ�I�����Ea_�y@;0,���3704�R�I�)�6k�=r�H�����^���ʠ�}W�����ϼ}�|�~L$K���=�ަɧ�v�yOw?�b88D�+�]f��	wj�s�6��g�䉖2�4��v�g_�m��i�^z���lP;y�}D��AF�?����L���I�-�0�I���I��,����{�����'�r!��C9�9\(���������S���6���0xB�t�E�$�*��?R5s�����+�} �G��!�Ҡ$#��H	�4���:4�s���Ic]�w�����>C����T�{�L��ES��N����n�U�A|r[Mm!*��� "#kߤ�f��@' 1�h�N{ы^�D��q��I��Aȶ³���=�D�1��Þ�d�D+�ko��-��&��{���	�j�����[��@`Ew���<����&�sS���]�ў}��8\p[Y{�,Ac���pX���h�Ae<���$�)�Ms/�w}���|�z�t&����N�2��Z�W&�7"��7������2���#�
j���1K*����q�/����>w�ҍ���f�o����򐧞&�9��呲5���a��ݞ�-�Qbu��d�4����aʁ���W�b+�'��0�Bd��!���NW�p�ͼc V&�:��Ƚ�T���+!�+	i2��M�7i6��& �5/{ُ{��/�K����9��D"f�䨨bދwRn����e<���K;����L���@��y�ޘc4i�t�w7�|��^S�"K�Y�xўpYe� ��V�P�n�&��Ǳ��C��N6��7�4�3� zu(��EQ�S�KEzt&5\�.��pv��m��aۅ1���^j�X"-ƥr�:W4i`��#���8�,� �A�R�u(!�xSc���_�i&E�=����OїZ���Ķ���V-,8,�CN+���?0�v���61J����*����r6[mXeh�#=Z0W��!�O����$:`y~�w�c+��%ɚ�a
@H��4���"�\)8x� �@���K��O���k�%sL ���X��r��; �MP��e��zJJG��i gA�!���`H�e�8;Fd�A�af�*��@3>�x�≫!^&bN41<s�ԯ�q�T�L�H�H�w��6�w@r0!k���f�5<�5��9Zo���-�
�G�O*��N��bVr�;��/ =@¿��!��5�U��Ԑ`���eƤoT͚<r��AraU�G���i�9?7��[�5�Z$���,��&�E6&�����71��Z��KsHQ1�Ԁ�w�N��\�4��Eӄ��Uׁ�MU���׏B��Y�$�b�z0@��B��b�i���F�-�t�fl�+y5k$�����m���?$��Mws�C��P�š�<����Y��Ɔ����Dh	U�H�X�6Ұ\;S��á�� �a�PA&��5�\�/��H�&pp�Va�;��&� =�@�C�\!Ykp��q��t	؂a �cc W�p���
��3n ps�*��H����0R/'EKRO��@����(݅��T:�9H�0 4$�|��(���YW���,�3<�����K��K]�����ye�06�S��-�CVnm���eײ����92� ��w�C�D@��`E�Z���4�V�Z�l4�*�B-V�Z{7��%�C���=)�]�iHJn(�Q���b� }���L{�@/�?��̘����B#]2�I�,$?lj����	��V�d
o�A`+5A� $�B�� �Ky��c���������I/a�h0B�ɓ��Q�j�l���p!��Ea੯�a4�t�Cͼ@�8�B�P1�H�|�DL��%�mAϒ7�pr��J���c�C���5���x�,$y�m��)���˚DF��cj���H�z ��a,<�Ƹa J�3n�@�8���������9t�'�PAY^���L����B���鏌��v!��k��3֒q�n�
?�Z�y��~��{�\�ϐא�ni����\���{�%�w��J%h;���fg�:׫n�o7��ɝ�';\�nS���$Vp�tzv�Ƃ����Z���H���9̛9��ʜ#����#��,F HL�Zڀ�f�����9�Ym0�r��'�+�<j" *l���o�SŽ9Dlt&�Ŕ���i������jZ��e��C��x�V~F>��}7�a���Lu5�yK|c��#H0�?1iw����34H��`��[��uO%��AG�aH��n8�*�1f�_�-e?_�P�KJ����I�$Bļ*���QZר�[,��3��He��3�+Y�=� �\AT�tǵ��+�>�LM{G��$P�lْ��!�K��Bc~�b�\��()]j�e~蟼E$}
����?0�UQ"�0�sn4.�$� �??����ĝۋ�Z�<����-��� �չ@��묭�,���I�d`rp�f݆��ꗿ2{j_� I�!`�8��k9��R4.Bb3ќ��d�Sռ�`���{f�G�ќ�a���[{��:��I��9�I�b�J�g��CF����F��<0��a���`�fa�	 {���������\�ؖ3և�Ƽ�h����?{�f�7H��M�XS�X�-7���D|�FX�E\�R%;l»M��tjD��|�N��N��4ikj�!M4i�b���I����jj��ׄN�����r��@�"�)!@Wq	�%���(��Ɯ�A��T�L=���IS4{R(?\#_��&�K�&C�[���	�2�,ͷ�M*!��6�[g��M�[�k[��0ng���:�����nrJ��sh8F�N!�=���oe��,�FsL��/�˺p���4ڏ�'R�'�'"��aR���h\��	D�'Xyuq+����˳D���W��Ը(i^�&��Y8�dAA��K���z�-h����>6���06�,��Fk�I��(mR�4Y�]<I�������֞�&	P�H�B�V1K_O�C?MN&)[D��P����B���AjH�O�����.��#@�Z�`�(I_k/��ԅ/��Dr"�i!�t�(�X�g���'iB��S��i��ԦEK������(���X��7�nh.��Rv1}���GK���k �Sg�]����:�ߞ�����/LZ����({-_�.�HZ��3����u�x �/�F|y&���H�hz|Ƴ��F�?��/�$ոE�?|MB��v�����9i�8jRW�I_����_���S�/�ik���[�x��a��3��2�B��B��$���.�"�"_�^WO=�	R�߮�g��`v�У�n�X.��P;�G0~�ż�f����Ŋ{3t�����7�I+��+C�6t��_�Մ��`��萪�ZJ�0��'�OR���Ii),�Fh�����Z ��/%������Hת����;D�b�2슩H��~�@�WذRM�=o�j�� &�k��X;�W z)Õ�"Mn���z�W�DsǵbLi��U�?��_���q9+�<�y��(N�K6>6n��l��yf$;�����ؖh���B���~���C��Ԙ�6H�b�i�.�#��g�g�|Ye�䩛}�Q�����~d��ضc�×##�~�/<�<7��ц�GiH�l;�?zj���	����\eC��9j�>b���ȑ�~�l��9g���=�<zȞ���|�6m�h�~֕��#�2	i�+Y)e��$ &�jË��0�"�b��9�d\��6�o>p{x���i}>�w�˹�<(� ���&K�6��8��_(/!N��K������P�T�m�<�f�K���a���n
��H5�� �.Hc�Y?-I�i��R�R�MR�$i��\wS5=u�L��Ik��9�qN��pa�?f#�9���I$<��w'�@Fa>���g��51�T�*¥yW_Rƥ>�{-Ո�YZ�MPRz����ƹ��J�.���K]>�V7�g�1K�;�-����5:uZeO��Yϵ�G�λ�2�Xw���C6;��e!�;^��
�B���L-�e�i�]�����3�58�����k����s\�����l�Ęu5[�9j߹�[v��~�֎#�7�ȁ��/�/�؞qųm�:k���b/��푽�����,��k�z�&��)��6W�q�.�;�l>�4��O���A;��>.��/���E
%/�p��\�����䬽����D�MN� �]�4G���#.g���(ˮ����x(8ԑ=l�tf�ds�{��o�|�0���f��E|�>Ҵ���#�b�"Rq��FUե6O�KR��G�<�h�B�4��u��_�/Ҕ\H$(��K��Yi)Ϡ����������R9+�Mڀ$s��&�$+�O�	6⹂I$aӔb��� ���������jIpW�N�R!���|�[����J����y���H̓a[���{ ��%���>i�cr<y��E۹�L��-�Çp}��8��`�4B]C�Ƙf�u���'Б'l$���h��q.0nn�a_��ce��_��b��3�+��qx!ur�l#˷��笿��s�*��>��O�5���o�T�u�u����!܁H	a�ڴ��i�z���s׹��<W8j�I��,�^�L�">��J��2�;���Zm��mނ�����unԍ�����OHvP��E��q��4�4�Ţ��;%)�9�fg�!w5<E��sK0^1=S^Tb<o+2l����;����Ѓ�
ߖd)"L���EA�~ˀ�7.�"����~� �ȷ|�!�#C�+�I�`=1 =���q�$6�+��1>b��3�m��o^��)����>o�L����5������	�AzG���uAӃ%K�h�i��3�3�^"���=��^O�G�A�/A�<Y��|�#]�N��-�N�f?���m��u�ٵ�Lв��/"���f�Uw�}����|N��p>�v����bXp_R�nX�6��V��x}�ݻ�m۟�tr�o
WG�=���5[Hw@ �ݜ1|�(	S�n��'�	~+sd/,Ե�|�E^.!}�=ca��0E}���u�~/�⣶������)��.�E#�	��I�٧��޷z=z��SY�p��ށ��@<�ʔ �CH�^�c=nsS,Y�А�R"���W� I�J�,���u#*�\?xa�Q
!�������1����<�f5�?aZ�/V2��� ��q�He�Nޖ�] i�g{��Q��w=9y�6�=y|�M����]�S@w\�O��د��hIr��@�8q%ozӛ|O����M���<�|i����q�w�=g�����졠���]�r�ssպ>r0��z���n\>s�9�o�#�|�=Y���'��N?�f��2�r���b����8a���I� X�����{��zo
�0(=�`.:v�d�=��!'`"n2���4�}"ps-�0�`�>�'�=��s��.�;$q|�\��绑�MWg!X4�#�+R�W!"���!�6�5sĿS<Y�3��P�]����w��`�0r��
��DF^?�����(jᤂ�dw�yH�Ja�A�O],ӄmJ�,����0��]��.�=�iH��M N�ϞZ��f�����r'eS2�e�9�	:_�e{��R5סCm|�~�Xs���(�C�I�x)�d�3Ns;�Ȱ��FAc��_��bm)��w�w]��z��9���g���Ja�y?ϣ#Ѱ\,��~᷂�d���*u�M�l&'<��bXu�
~hk8E���;��[�}�1�Ot�_����Q�[Bɯ$�B����`?s��h�	:IS</ۂ;��Ç�ك��t��@�5N�8!aa��!%����	���$���6��A�<Wf��8Q�[���-�Ik(��B�?��9��t�P����w�RE��P�,�ʮ�g�k�sY��V��!���Agh\��܋�QV��TZ��#��
��&�,6#��;�+�:��AG�ĖD0�]m���ޘ"�~i\u�J���hrm:m�6l���-��~܎�[Z�C���Zr.Xs��C?��:�m�v���\�p{b;�Y�Z�Y"�������:�>��KS�$�H@Nx�?��oL=�rcn�ȿv�v�8�-��f;H�%O�q�~ѓ��\�ŒQ��@-<��o��ou��J�KCB������!*¥�tzϲ-||�}�����+��E��|���/G/�����5E�Bx�f	6.��K�5��1�L��eRq���H�8��Ԡ)b+)�)H�g �@�!��I�yF*&���i�J�8�gTq$h���;c�u
xR�0�,���H{~Aw�;�Q�
B���֑����P�{i��5�N����6�.��'"?��/��~p����k����Ş����u�ξ�w<���۴%F���!������Ǻ@q�{o>h���{�j׭�����S�8����v�#!)���I����F��w����"J��+��:� ��D8�f��Co�Tq�=w��u�z�>���G�p�d�+��6�7����x�8:fa8~֯[k���7o���K�F�8V�z1�R �հ �� /��W�7>�r���� @`��$aJcL��]s��@1ȋԽkm��VµsΚ�fPU+8���2��-Rz�W(u7��`����FcG�A^;���.An�nƌZL���%Ė�����3]b+��&��|� �fL�l��́�3?s�����/^�,cQ�p
��{��Fڀ$��(\��U ���F7<+'�b������3`>Ur�4({��}��r�o�]NPx?������-��|�=���yO�V.U\3��)e�UlR��m!J���ƥ6Jҭ���3
sj��?��n}d�|~�W�ӳ UR�Qğ�E���i�mvg�����u�L�>:T.����mf�������W�ǟ��Uts	�|;�XȾl���0[A���^v�Ka���?�G����	�kQ�B�휟�)�oF�8j���~�E@U��<M d+�X�y�>ג�� H�l�~�n\�@4��~�Xx_���ᣨr����v�H�}���E�\�A�07u�٣�"0�b&�#�0>4��۶�w���a"S%������{đ��q�wv�k����`��,�0����������x�5�$E��������geQ�%�#��<ii���)��3`vc�+̃&�/5?�J� ��!M��������@a�	w�v�=D���`�����e�4�ǿ!H�!�[���"R�1�A�|�(v�2�p��}�=7*j/�-�	-���H��@���y�!���:���hI�'�e}��7��6�=�-���z�LO�ځ'{�#y��y��a	
��=��0��[�U��<B>4b+���B���x�A�ǎ�5Q�9g���89;r8�yb|�7.�g�{�My,���@_���F2Z���	۾�b����c��[��={
svȃ6{[��<i#|�U�� _�ڇ�Py�]��gن��mnv��ز�n?x�8=0���䙢��u�]yՋ|s�H,"��� j x0đM�	�x��?di1x�Æ������TPM�?}4�&�B=H9��7!D#��0�:!�kæ�c%�l�����@�k�l��aO$��Ę\-��9�Jf��a`���^Z�$ߴ@����:�%��7}�N ���b�� d;�w�G���CCX$� -�F^Z���y䅣��`�ߺ¯��n	����A+��F)�~C(0C@�
�/�q��ay.̅��YCT�O����uF��؉2YMa�J��ܰU��)b�zr-�C���E����>go�h<�a��/�@�U�����!�̟� ���P�<�g�NU�V׎]�b1��|5��#AZ�gsӁ ����
w�Q�+K��o�F�2B�Π;��+�)�N	A(c��p�Q�,F�<���)[�R�P_������oۺ+KwrȎNO�����OJ��9��߲y����/��Ns�$���vXj9��v��܀���5��l�����e��l��.xz؈�@?�X �U���۶�U�}�o�ѱxp�q�-`�&iR
�#i��?b�㏹��(V`p������!�'�?�CA�ǵ4l�|ۍH�Vؼ�J �@���ߍ, ��-w_��yA���ɼra�b����Z�x��H�lP�~`.儗�(�g��"� ����9$�)I�)���T��I�o�&8���AH���3���'��a�;�d�L��W-����@Z�����u�J&�� �E����7@��?��%Mr��~��k��� ��?����!���3�:0��"Θ ^0�MK�씌�uG�e�L�RV3/�a�d+e@U<wU����|�}����"G�ћ�^w�u��[�Rd���0ƶvݨ5֌�qT���[��� ���5�܂s�p>��͠C�3������y�u&��'��[�/����#�$�}���+���Mm�94g��k��=j��DOd�ư��watj8��h+���w��[Bɓm'<�Ԕ7}��	/�@�<O�����>������7�����U��x�Y�����-��@ H8<O�B��<3��g+��"�Lĵl$
�R:�Z���5ힻo�COl��Բf#fW���G����׾�]�<Z�T�20����Ԅq*~�"z�c	BB2�o�)/D7�Ad��H��F�5N��HT�$E��Y*j!��4Kg
�(��pPyh`���� /��#El*�k��͡
d�J����GՉ����>���9hE������"B$d� ��{�k ����_��B����a�XO�-��3�
�u0vy.)/3~��++�F�f��"L�70���Zs��G� 2����'�����=�;��,���y�� �ӷ˯x��>���֊R�ds�A����6;�̈V�W�U+�%y#{��d�>�����^��Z�����l;���W<�r+W
����gO��2���{l��=���;β��0�s66�ƾ��o���E���&�_��I[�:���Zu�֎G�M^�z�i_��F��Q鐺0����x��Ojz)l�@H<�Z�y���`S(=C��G��`q_n�]�u�ɥdU��k������ᾩ���Q�)�V5F4�[��3|�˓��≯�����UP�M�S�����T�����Vau�9)���)���q�D"T�C��	���i?��-��`R���ai��Ռ?����>�p�yS9l���i���^�g�p{�rL��F�V��)g�4D�[j[`�� %K+Ax���)�.Ps���N�����ξD�C���Ʌ�w ��H(������.���<��"s��!ӟ�Tu-���H�vl9h	��%Z�iI�?��ʖpO�3Ʒ��Q�Wݏ>��(�@8K�h�/�>�-�~#��I��<�e��W����0���w��{~���s��;�|�^b� �0g��@|��p>�v�eW��݀A��@?#���/}���_ז�P�����-�S�ֺ�폎�I���l^6�E]l�u��9;K Ҽcmn$�t\��$k>C��lⷿ����t����jc�[���o ���d�%��qVZ$�`�c65��L!+��-0���{0x��y2�h��-���k�Xz���p�qGc3C�f����Z��	���F�����!L���<@`�/�\�t_�B(���hi}U1gɨ�ajt_v�d>�V�z��`��Щ�������ijo�zB ���M�M\X3c��)����x��|x���<����%h�w �5�ɳ?��O!`���{�����+�3�:ׁ�C�!�h�q��ٻhPt��|�рphh�|�f���rb��>���_�^D�	��D�zZ�|����<p�9d��4�ݤ~���.�S�}C�!!��J���0��/p)��$���������|��a����_���-�ܵ��5�����2`Y�J|p�}#st )h5c�1���������h��:����7?_��x�v?��}�߿�v|d43�M��$��O]���N�����	���#	pPq9�GZ��_x���� y�J�ݖ���_�5,"y����A�}r�3�T6���_�MsU��[�!�܀- 	��i$�N��,��=�q8D^:H�H�ܧ���ڇ/djoJ,i�Xq��P�t�P5�����9������,����RJ����
�������b���]���d��F�	?��s�q/*���9���n�!���ј�Ӂ�	��0�o}�[�>��@�T���@$��e�<���<�Ϙ3�@��<%~|��0����m�>���o���<�,T�JB �g��Ә+�=�va\.�7��wF�^��=" բ<�A=H���Ʒ�F��uߧ}�Z��@P�]F�1v��_�_��~����(@�g�g�D}RT��cM����;�~Ͼ��[��`�w�3�y�B�A�~؞x��� ��'��rWЅ���C�?����QJb�:����&�`�>�s���\�&G�T�M��o��$d�H��ˠ�$��H�HLHe
�`��y(+d7�K�0�з�vچM6;w8�;���Tp[>���+�,y�k���^��(�'_~�����W�jw��N'���d�|���$?�Y�zQ��?�;�`��.UJJ�f���V�y?X5�1��H�iV��I+��@0ހ�0��� �!�z�_�NEf��yF��i Ҵ�r&�њ~\���\p7�̃�} n�� 8,NhG��U^�����}�<,���F̃
��{���T��Y�����_Q�i-
e>�[���
�×�I��{�5i�*��r�`�%A^*���%L]X�ny��9��zιچ����ѽ�������-�:.,�m�M�؍??�`�\���GJ�C�Ё!���M8�gl$�RΆ��8 ��R��F.�^�crk�0�'���}Z��s�V�\I��v⛷�!*`�<�l�NW"���A�'��z���| ³�9{�k_c?��{�U�q5�|!��L��Ar�4��ԋc8vQB�{�"�JC�q۸aKP'��X<&9���k�{)Q��د F�=�2��G�w�t8�O��?��/��s����{�<���v?�ֽ�E��?j\~�3��P�E?�B�^�Cب$0Ta0i���A��N{�e9)4�t�s��t�0�2�ʯ?��&��'���^{�΄xv���(+k~���p~������u׸0	��+Ulnf֦'��?�
������;��soz�y���/{�;��5���R�.����4׿`(E��9�ŰR��bR~����Zנ9CH#������,;m'�B�K]S)Y��|�����sA�:g��߸�=|:n(�sO퉖��6 GyF�0Tj�Ԣ(�Ja���c�q���ȜH{!y�sWo��`��sG:Y_�8��u�s�棞\�n#h�=+)�<�*|'<��*��R�ۖ�< ��7�������"�}�tM"@��#��
��:��Kv�X���Ar��q������"щͥ�h@jogѦ�7M!�R� B���1�~�����ʴ	�La�O����Z�]Z�\�
&�'D���P����*�U�&L����	J�z ��|8���Z�x"��5�,�f@���ۉ�	GNSU�,$z�w\f��q�N���;I�����g�����M� ~r7A>9;�{����TԆ�����B�Q��%,��[��'h��k���b��ҡ�\�RB�+t�#M�j�
ԔP�����۹��.�b��9U�}�������mQZY�EF4{���#������w��!�w`�$UEH䝣w,�:64��
�p���t�q������L���=�W�L�`؃>C� ���z`��4ߗ�+0�Ft,FDy�H2^v~���]�ΡZ+7��g�k"�\�;6����3��#��3������F��)"��n<�u�!aT��S6��
b�Y�<0"�C%gx9D^�00
�h>��3�A��Nޖ�ow��T�b�� �i5�iz"����l|�tX�u�+�=yȓK�&��z�U�.$)�Cl��[,��ڮ~�����+p>	i��5���c��=��l/q��V�'�	_`I�;�x�V��p���\}�cӶb�u��!�$�S��S��I��x$�
�Z���_�B����=�Vn2|��+����O��r0s�T��SЄl$�z��?(& R�ŝ�.>�&����&���G}�:�$L|�B�f������O��HS+MAƋ�ϻa x~!$ +��\|��/�4}�7Z� o��峂E<15C4 �ߵ���m���)%J��R1�0̑�#Vܷ�6���6b#k�ݘ�̗��A������Gr�T!�ԾM�4��*���qg���V|�O���\�rZ�4�*�*q������+xBը�3/�(�5MӪ�J�<�n�������=V��
.�P6[��s80(��
̢m�����ʃ��̻K'�+�B$�~M����J�P�Ӡ���ru��M��V�&�=-+)�1~�S�{h�N*wG(�N~i�"����Q�$d��]i!t���1�g�����!�4 ŀ�]� Oa��y���7�_���o�t���N�Ȗĉ���j��ٓ�r�������u�6�E^�q�}�8B[����p�����mG�J��jZ�+x�����m��I�5�-��޶ԋD��K���t>$]��<$$��`���\"�z�H�0Vmn��~�d'�y9:L�8E�0$r��<_I��X��c-��@�d������=���2p��VjE4��DL!�Z.�YZ��\W���ؽG�f����!u�@�U�K_W���Y�HN���i�g0FEz��k��%�IWM>LHbh��0ϐ�41e,=բg4�Z���px�N���x5k��o�38bs�i/��C	E?�H���`m�s�s�+Pp�m�A���~�	R[M;�u\M<q%�+�E�_���(:+O�]>�*�-���I�4a������?���\ j�	+H�5��0��b;��t�d/��uJ��!��k�@��-��iv	P��ޗ������.3M��p�r$"t҆�Ҽ8+51NͯR�^pt�,��ȴ&����LS�5a��GYYaH$$�xs��"%����"�a�J��E_�R�UeA��Q%2�gb'o�jQݞ���A�G$.,���P{?�z0<�H�{)����T�+0����ƂI "Ÿ�|��Śq}�d���=j�� �!w�=�1��l�_����?7�����vq�*cq8#l�\ڌT�M��$�*Ǐ2=�Z�4F`%�*� -ō�v�el�dÕ��$���F���6�U83ӳAI
?��Ē��V�9%]��%b�������@ɾ!C�r�H�#�m#WB�C��[IЋ<md3P�v�B�Xk&�Hާ<@b ����$�9�v�
`�$e��+6D����������j��N�&AFn��ߒh�Å?<b��~g �5'ؕ�׿.�x����]�/_tXO��D��|�U�����,Ы�A{���D����K���^e��TX�=y��'�9�_�è2*|;����(����cc1hfzzƯ��"
u4���`Iz��O	�
�N�`~f��w/���$��m�}��wY�Q'l�V݉?Iܦ��V��(�V��%��2�����?{|V����� �:�҂䛾��%>�)��Y�J�����vi��
^i��C��u_��O����`���=���Dwzf�/xL�.5"�܄uMZ'���=�Y�s�r%�ڹX�qdl�|U�ȉU4��n��,PP,�S���i6cpY������������Ҧݽ��w$/��^ӑD���y�7�Ʃ@�d�	O�;�)�^��C<U���g�s�:�FFǭ�P�#A�{�὞��۾��݅k��H��+zR��P4)yO�Y�������U¦��29{#��byh�3��N7챃�V]h�T�(��V�+���]iW�טSb�B9��k��Ȩz��jO��ǟ}��J7�,I<�j 6��Mw�P���oqfn��5�]��O��aÒg�`��H�7�C&c�����Od�cCn�y�[~���B�]8�k\�)��'�
���ύ����$���B��֬�Ds3s���cl20����ƀ=i���N�d-�2�	?�Ǘ�>
?;�>�xW��S�n�/��]~�v��A���K�/���4��
]����`�dt�_\�E���na�Hl�tNۢ��i[�U\�y�G�N���U����;<56���1�!5�۱�Ѡ����)��j+����S�O�w��%ҔN-O�'���Y�EϋB���Yg���m۶%�Ջ���!��9'�F'0�3�\:<kÕ	�K��+�3�,�w�K�/�}�C��L�#��!�I���{�� ��fi��3�lu�����);K��k�(4;�o���Z����j����)[����� �/��\��>�����]#l�:���h�T)Lz�"��ٺ��ڦ�6xpɸ���|%���7�t�둵��E��"�*�n�N3t���C�BP]�^l&o��ݲѱ���uWu�T�fe��"�?}ih��(<<M� ����+��jA[��O��o�|��%�L�����\��᜔����yخC�q�����G&�����\��0⮝Ĳ���l
�D��Q i�3M]�r�'�}�G�񩐓\}_��W�}dk-�"�E�!��l�zz`L[����rm$©O~�N|�?��@6D{��?a�#�dW��S;�������q�0p�g=�6>����Nد���{��'WA��{��^_�`7�s�N��_�e�5'E .}^�7�@HS���FU-@�Hi6h%*�%����s �'�-�������0���I�"���*F���T�[s����ک֧-c ���O�<V�˓�$\�-x����CONNۚ��6::�I�<-J�-����b��b������zh��>�������)�&�lg��L��5��}s8�s6��}{w{j��{���wv����3�+v�gۛ��3�����T��z����G+���2�F)}̉�m�= �nn�ff��;��O��������;�ܽ�v�=v��/�ˮx�5k��!���h�#�l�$�"������?��/�c`�t#K����]��g���v;p`�x|�MO�Y��iFEIڎ���A��p|i 2<���(�S�	JS��%���}��j����	�G�,d���o�6q��������z�*��@X�٥�=�ʕ1��j�A���Hު�Bb�����E�%����vw��l7�3?�3.����ܛ���%/y��:�L��$�i�����曾���,�p�n��[�v�z���v�}�:u���կy�}�3�q&4T����}�|;yO\���K.��Nߴ)l8q��s�MO��O�6O�7��2f����_��?8m��ɟv�<�iH�7�LyB��_�Wx`�?��?9�ă�҂TA��y�ۋPJ��߅Џ����n#;Ƭ�+[c�aL/<ݦ�o��Ҍg>̼Iq�����2�k-����ׯ_�M�G�ŵQ�g���?ӌ���_m5�S�T[�en�� ���'���ݠ�E[0'�F1�jں��v�E�:�Ǹ[,��-[�Q�
-e�(s]�`�5C,I	��N������&ug?F�׺g��/�T<+מ�C�=���vn����v�Y>�n�_��z�|�]��gYex��=w��w�9��[o?��;�ߖ�eY�� �w�9�������~sP�6�y�������q��yN�`�n���l���<����Co��%������~��=Ϸj��+H8���˗���rVϼ���#�i�U�]��:Y�x��+x7X��Wng���Ă��O���al�K��O����P����D�"����$#li�k=�T;Վ��׿��;��<���h�b.���7�5�ގiN��6��;�!Y��?����:��I����|�����{��p/��~�4�=��kҝ�|�@�����پ}{=�y�w���G\��ʗ�����}Ǩ?w׎3��;�<��;��?�C}� �E�۹ABŐK��G�c�6���[�G�]Dܻ���1�H��qr�?��+|s\p����o��B�F*öo�#�W��'�#��^|O���U2���}���X�QQgG�qQ����;X��X���y<��@L~�B���/��W���7n<� x#�g���t��RGS��ޜ�P�R��Ơ�S�Q�������)���U�:Ћ�NS���R�S��K�'_Fp�U�ߧe(�q=�+`KcS�ԗt܊9�8U4F��\i_���VAy	i���K���{�0�]1��$�-E�g�]o�]_���!M�R<���)�{����x�����FYG�N8�`���-Y��F��~���'7jYs��~ʮ��s����w<�~�g��fP����
��D֭Y�$�y��]�ن��lٲ&m�6_������7�j�-�����i���V�Pz�}c�\�R�tϯ���Ŀo�K0~��o��a��}��y��m[��������n;q!��������o��o��s�d���q�ڵ���N?ɿ��� -Tgڡ#���U2�p�dxdµ�4�9�L�D�Q�����PM�1���o�#��}���چ��tɪeL�)��C_S�_DB�S��X��mpe=��V��-ՙ[��{�oH@EXD��h]I�����ا�`s�*�w
��whR���+�9H�$���`9�+�\I�y�{�1��d��4��]j��zi�)Q!s Ƣ@4�W���[�S�I�и�GR�b�$��3�-%|-�豸�Z�1�l7ݦ�Y۰q��E���	`�;G��ƈ���6]�-����� �R���zd}���&����w�<��mXw�{��fBok.���M/�[ȕ�H�=w�m?��W{��*�Ɲ�w�b�y��v��N�d����XU�K�e�����AL�Ng)��г}�ͫ��!��0���P�|����M7�@�\��?�zB�c[t�l���=67�f��#G��<'���I7�E͉<�}�o�o~����ZǦ��m�HSɑ�BL(F�}�V{�������	�KlzpP��L*��L�k��"h�LQV��T�Y�.�g�E]��p�&���̝b,��k*ً���J��q�͈HZL��k|�Li&iD/M�O�h����x��� A�&02��5��B�T�Q��<VR/�TkH�N��1����7Xn� j@����h��5_Ms���'gё�Dl��}b�<R>SWg��᣶���m<:��5�Ǖ�
�7�%Y��esl,F��x�nإl#�?s����^�B�LL^9�8<S	���Ӏ�����`Lh8DB� p"dAspG'�"Li�R�r�'��e�(lT�c�ר7|qt�I��l��hZ,��TԴ�js�Te���{���[n����]WP���fQ�vO��g-��ZN����:��)T����(�ry��<L̉���� /$�|��y����H��d."N_qW}����Z�n��!���<� $�RB��M	�E8���ko*���I��N��4'��X�����ԝ&RK�r�W�%MC�!e
),���1�=�\��z�l�E�b�������� $'f��	��>����^�֐��]bip��A�RoTAEiiG�=e�;�:M�N~Xiv�V�]5�o���/�|�ݓR�M�W���B��ֽP{܏e���ZexT��4/���+?��#�#�c��9J���p~p�云�1��83�%�R#�Sw�6O1!M
B�u��9.��lxP��'��i�R�#�:b��G\Z����uu1HC�l�m$�[��Vk̅��݃�f�N�L ��}�s~ )��я~ԋt �����A��v�o*6�b��Z�0�9�	kRM)l�E�6O`R��3����,�v����Z���~�C�f!ց������)/�ą��`�}I׸Ѧi-B"����酂t����m��B4Io�1����N�s%�J*�4-b&��S%u����MꛘIJt�0oiM��_f�#�Ҷ`+����]�D�G�$~ER;�'�j 
*�I���<(��>�K学��Ms &�{5#����2�*�Ij[-��\��z\n�|��*�z�o3�?Vm���p���̡D���I�@/�������Jս�0���g��?�^���\;�0w����m:}K���@V����"i�7n8�?ɮ���c���K�4�{�C�	O����(�b�*�/�����a��g���a7���xҬ	� 'ok�֨�C�<b��[�T�3t�Dx��Xt<f��Q��~ac���\:TIWS��h��S��d±�y�c�
�]��6��Q�cY�T�f3��ii���`��}�K_r/ ��W��U����&�w�Pe����J�]�����T�?H��6R���C��ߒ��{H�ZYkŜ+�j�7ˈ*$�H嚛�r3����G�eҤz%��1N�2'1�h���~�.�`���UW]խ��/����uBJ�L�((�)�EED^k'����:i.S��bAz�$5�ߩ�Ͽy�~`��I���٠��-�l�t+�Dx��O�.E���ͯyJgR?��x�N;��	;p�q_?�w�w�%�������1�o}�[. ���o�׽�u��4^i���K/��|��#���5�"��g�T�u�6;�z�ӂ���iB�/��밖-ըV�Nx�?����k�,xp��]jc#�b�G��l�c�mzf���IĂ���Gm���v����!����&�j��w��~�w~� �R6��H[06� ))�F�֢�I�g�B;��KʡO������!��Q�����a�b�v���p����GV�č����
cÞ��s�׀�$127�Œ��\�P��Qaih|ǵ�G��Ԉ��#|]7���o�%�{!xz��J����E?d���r�|=�S�O�+���`v��u��������������g0~��7��>I���h(���d/�� �J|Ιgx�D���%H�h�A�i�,A]���>BK
ӉQ��@�觠4�*R�+���;�Rږ<���է�^�Do��p:��"G���O[����'�l8��k��f3��2�g��U�f\Pr�𑊯K�:���^W�o9�1����Z�?4 #����m����{�Vu�"��g:���6w���5�,�5���k��Bb'>��dtc"!ި��}�s,$��7o��[ny"0���P��DKk���?�.}Ƴl۶���1(P�߯l lr�5�4��<h���җ��Ŕ��2$��C��������=?d�F�8�p�5'���Ӟt�8�� �>�|�x"�M0n�'��D�&����F�ĀM�
��� �,�k9�h<HFƆ&�!๤��`2_�.���H��@8a��%!�-�l��!A���]|�Ů�+�"̞���w뭷v��@�!>0<�R�qE�h�It4�����A�!�`�3sG?��O/��wa8�^�>�����b#���@���x�'�42?ϔ��{��W�H柹�H�x L|Ƽ���\�#&s��A�b��ꓰ�ZJS�N�0w��&I?�S��A�EO��Ko�f���!.j�x��pK-��?g�N�jW\~i83hay�T�ߛ�eU2�ļ����3c2pb4�����e��A�0Rh�'���a��O��w��q�96_mط��M;x�q����Ex��v�%�k��,n�Z�;�;��^O�r<e^Nx�?����G������U��~����g_ye��Sv��ٶg�#{�ə�y��~#\x���áYX�S����1|��_����.���ȒhW6��5�yM�����Յ�-�����;ǼH�R!˴i��G�.�wo���^0�Xp:Q*,"� !�^�
c��"������5�saTC�s��0��I�A��������"9qX�~�p��< ��%X66`'y� ������Յhn�
qހ���?��3gR��ŕ��<�	.��ox�"am �H��ƚ2<��t\��[�������#���1?�@<��y6��y�X��w�ß�e�!в� �0�J+��z����H?���v���B�w�O�k�����ؙDj��Q�`r����=��nl0"����#�´��5�����9F�Zj�Z�	`�3`���;��EO;;G՘��J�8{��N��w�+~�5��.��מ�c&����?��.�ǚ�ߘOՕ�f�\��0`���c����]g�sٱ.���m:�p�+�a��kk�m�����H�n��˩
:��ۊg�N򖺖�0H]_���H
�2T�3w�gO��{�F٨�����t�MN(�"/!#��g>��@��90��]����)L��r�pl�E�ߴ�Pζ����*�@���ߎ�����+�(>$���VaqK��vߧ���o��*t�&O���
�8C��$^��A��;�⁔L�(BdyLAFK�ć�a <��z�R��?���l���BX����ε<��5��v��F��Y#�0DBȻ �Kpu8D���BZG��`\ya<���0��������\3��O�`2�����D��HPP�l*�Ë��H��^�җz?���Aq�����{�0�fO��y.�/���ó���jg^�/�m�� `�E����Fgh��"L��+���6�����Y�����A󥆯kP�6�`tl��ȯ7�\�/ʈ�%{��Tm�V�9?�N8t��Y�.�I^Br��������������~�;cK�N��g�3�v��}��b�]�%g���Z����O���1�+�aܴ�Ȑ=��>����j߻�6{ы^�O��G��9�g�a��c7�tC8��,I� ���w��UY�j��s?�sV��!�*�� ��QX�b�= A}��a�MR�uLK�(����V���A��s��˭��ѱ�OYA�ѹ�)o��֬�����F�5}R>s!� �8Iud����XUm�[Pb�D	�n��B�!��`y�C�3!�H�D'C����P"�qߣ���2�;#�N����!�2�)]8G:r���C��L߸��>�9�&3�0J�DzN��p�Xb���s��	�M�%�^�s�0�7�=�C������ɷ_�s�b�g<���	k�>��^<�x/ϓ��o�2��I�	�b�0��K��cXZA������vػ���;h�A�m Q�2b?���zw��w�c4�GZʾܰ!B{�G�7�}��Ky96�x��}�S��=�G^`�}�U~��:� ��e�Ұ�����/	�Ď19=h�Hē��q��A_��t0٬D����|SOL�q)��٨���Y��h2�	��|��ԧ>�Ź9���/����!X�WR�F[�7�����4f\M�b��P�e��@�[C/�\?Nl�O��6���B�|持��Ƈ�-�1C�������i�E�Q��q�H� �����ġ��sИ7��?�Y;�c�c.!�<�����!yq8a
4�H?�Fy'k!�O~+�C���x��$�2E`ƉF�{H�"��i�f �<�>\{��A���5h��E�1a'A��11�J���0*ր~ ��,	$"<�*#3sGc��H���a ����z a�AE0C��z�C�!�\#{�y&��z3_�����1�^�g���y�1��D�4��=���RD�S����΃�8;�By��]=��X7[� Ͻg?�*_'�L��g�9��=	�O�T���xff�v����n����Ӄ���Y��F�<��Y\�"��flx��t9�?��~߳�D󲯔��=;�+�y���^��9{$��#�_t�i%s�Ң
ד�&F9n���F�!��� �>�tH叾옺x}�vl??�3�67e<t�>�ߋ��ƭ�A>k�"����i-Vي��ϟ ,I���!��������!�G��F�c�:$Y5{��$�#�qCp�	`�=ćk!�ZS�!}�A�a�H��%D�y���_����� �a]Xs�v �:�4�OZ	?@9����!&̌�A�!�"���7Z��A�Ȣ%HC�9���� 0�����|���<m�Ly70�"M�^��k!��+���yd 8�Q%�A��}%+c��,����� ��|�o��~c,�V�j$�Ѱ�ܧ=���4�����4z/ۘe��y���u�].���gنM۬2<�I�b/#�gj��+:=2�| ��q��o��k{�A�!�1��)F�zMI��~�)�`����>�/0�=Q;�d���5������(�,Wm~n�\�s''��t�B��j1���/���
G��� wN��������Un_<��a�(�9_@9����u��D���kn��X��H2T��Ѣ�]�ɦ�v�7﹉���7<,�#�Qp���6z��J�Æ�@@88�D��o���Ɗ��R~��4\;-�.�7wfȔ߹����bǏ�R}����ɯ^��I��=H�rߤ��4�X;�ʡ�����s���> �L��&O��B�e`�/�[�ϣ�a�`��H��	s���p�>6�'����8`H�M��ɘ��O���y�x7��0�`5/�$�����\9�3Ew+e����@�����r>�qu��b���bzs~
���s�-�	����
�w=_�s�G;����ԟ
C��>���0/֗�����U��4'y��Cl�!ڂvkC�[���ͷ;�w;��ʼ�|v;���saP!X$r�,�c�Ĺ��&o�}���R	�$|�vb�W�h�4F�_��_�_��_w�3�� )�.�_wBɁH7��4���6:��B��!�p<���hƒ/e�7�"�|���4�q�����%��0u$�P!6V$b�{�l<gy���&�<宙F��^�S������C� ~��ȍPy��8$qy��7����lt��o���~����l<1�5�
L#�%	�@*��TiO��f>%,C"?�ٲ�X#��wA�h�B#A����G3�Y�xJK�z�4!}��ZZ�����$Qk�5W\�����8�vC[��J{��-�xK���.��ՊkQ.���z�������u2�	�ŹG�VW���cǝ�9C b_)c�������,h%��w�P���S'��-���\�K�nl��|;$�%�˝r����+��.^��|�qCG8�������A--�Ghg��)
Q��7�#p�x�B��</���p�W�Y�%Q��W��8D��`�N&DCɺn��B$0�}�E��d3(7��i~������o�I{�{�c��G����R�$u�ͽ��T���b�NAW���{�*`2��s�/��*	Sp^%�:�|�HV%HS����yz�,W;��
�V`��1�*xP�RF������� $��Rp}�s���� �Zl`�@�D��adozӛ���4��3�O����f��I{�A^\#�V�z¨�c:�2�k��'��	��0V���}���|ݫv5�5'�@����S��BA9�b�.@i�n3Ȝ�3cD�~P�.�!Q�����A]��ix
�ت7�}���2�6�n�DD*�?��So;	��V*��({����B�|'���R�ͥ�\њ5��� ����z�U8$�T�����ẇ�k���~w��˳GH���E6�.�K"�px�T�:b��W��'�nY�`�R�s���L۝�H�TAD��0p{��{�ԩ�5�D�%M��Hʥɏ;M�JҊh)���4�l*zF��&��RI�&��&`CW��O>��VD����oi�`�A��-f��c�g�)��h��]ஊt�D����ް��w�>1=��T�M��2"��U��[�-%���_o�~n��-�)�c[��3�/0�@�9����p����~��ֶ�y��M�f{�c6ng�n3˻&�7�F3��U���� cFg1O�W��񮶃���张̢0E��R��e��CY!�N���2�b!~��V��ϧ�+�\�&��Ri�Z�Z�v.&�r�' ���B&M�,Ҍ�:"N�p�5��:�{�����?l䃇��Ƀ67{ت�S���RD�$��v��5,�)d�I[K���?�%�J��Y`�TAT����q���H�H����C��xC�O�囘� �x�=���E�щܐ�	���&?�7ݣ흤�D��/4lt|��v��*hxl�S:S�	�A��k�-�BSFtN��i�i���\�f@�C����w��#��Q𿛭�f�t�
O�v�$5�jC�Q"m�W��w`�O�V��b��XʱPT*��E�)%y��3('�6-5�*�w9�Qj�l��8���x��c�Xo�@�|� �/dϴ���$��9��)#'������ϵ��q�?��=1�����sI������~���o��0��1�H�T���[;&v˵�-aM�%f�g�=�����5/�a�Uv�}�&�gl�m�7F���kڙF�g�`K5i3�UE���������vF��Eo�J	���\����^�|�[�J���d� $��m��A����S�q@�C�OE�e����� -2��S�JM�y��;���}���{S�}+��V��sso��9�����k���n�bwio�ji�I߽�_�w{��٢!(�8� ���=�y�8�Ѳiy6A�u~�l1���g������ ���o�׎?ꖂ@�y��`o��2"�ԭ�x.\y�%>c�����,b�CS�y���t(�"xMj!�C���� ��$E��ԷS���(9�QMk4�b��?�JX(��F�.��U�U�<���^z1w�d7�HǆJq�w2H�c%k4���)�.#F���2{_5�q�8/�Kl��٠�F�c.�[�,�1�[��[¿���{r��{��l��7��1�胱��-���/|ZU�jH(*-3m�F��m.mBY|��ִ�����1���w���ش���5t2W�mgƎ>�@�1����x9W��C���p�F(���K=�۟�7��(J���=J�
�5��}�m����(�!C���H��t�8��B�^o��C�l�S'-�rm��6��=�l߁63�g:�X��ke���BZMk���a�-�6�e�f .5�[/W0���؍��>�Ϊ�1KY\����l��_w��h�:��V ��*^� �8b���.*}�LF
��C0��'UX�s�=ç9㔰P:C�i6\�ѩ�C���J���{�z7kh��K�t�ދGB��&�W �e#^�R)2��Gy�i@��c����<��o?RlyY)=�S)������x��V��xtσ֜���Y��#�{�68�4
��c�`��h��9�i4�jQ�ˣO��c���֑bX� L�3zx�B.�(���p]O��f�GP�L���)�8��ӛ���pH�Y J�І���u��q�6z����\8��H���=���<?o�*�k���$ɷF�:ַ��M�ۻ�����gN�sAX�mf�4�jA1�4(1}l��u��l���^<i�A�GDe��l�m��Yrɹ��+��t�b���S��!�I+!AB_�~���X�ݳx84ۊEu#�a�U�ޖ��.x4b��ʵv�78�?¿X�� \�ctXO]�fpl�Zq����e@�H?�W�ݣC�v����ڵ��l	�DؿȔ}���:~���QF��l)�xQf�g���w�7;�9�(���[��thb����@��P/FF�o�s���դ)r��W�RC�9�R`J�y�K�q���_�u�Ycf2X'eg�t�C�+�q߾�v��;���	+v+1w8�~�3T0Js�(FEX�mW�
������� T{0;?��� d�H��9)��;;��-�'Y�m��Mv�5��=��a�y�aC�5�޼�;�o�s]O�hw��ʷ��O��Wz-P�����W��I��~R�N�_��_w&�^�9�?ˮ��*۲ꐚW ǽ�p���;wy<�{��.���ډ3�+v���x<��z�>e��,�x���꫟f/�����#�7�b��N?A�5:u�t�F��M�(`-$ �!%�L 	w^G�� �����5���^¿ ^9i���A.�?iǚs*!�m,�ȩ��SA���S�D ���}���g
R������?�`8C�sJ�¡��-���6�*�v-�5�d�<=���`��V�����1���E?�9�I�����2kU8_��ʏ����W��X%��9n�	�Xj��߲ҕ���	�ѽWE�O1(UO�ޫHOך>�����T��Y=c���2�^�:lB/�b9X�e
9�� h�M�c�a�XS�x�b"����V���&$=��/���e=c����y���ʯ��i�c��q{�w�]�4z.�����0�i/Ɯ����aՒ]v�v�,�`�o�����OkI�EO�%�Y/��/K��i5���`�o��K^�"p"�v{����o���M���~����.��R[�f�5�mgy�RH�*Q� �P<7}�o�[�3h���^+�����"^�q�	�L}&,Jf�y��۴����=웶������8
����t���Z6"H�� ��Vo�TA�f�k�8m�"�Q	c�$�T���u�W�Jx��ƙ/sRe�)ǉy�Ŝo�!���L\Li1��sD�s�񚠕4Q@<>\�^^�x~�)#Jկ���� .C�E��1�7�4����ž��(w��n�����7��Iqn4fmr�v�jC��-Y
mv;�,ve�k�f�s�&����f�n�F�4�������3�8�c�%;�԰��:���S'�ѕg
/���p���k�pf ք�si"��9j�zw(w�;lF�ú5k�&��z���Лv����W�h���u;~���DXl�w�];�ˮ�:�k79.�u�۱#G�?!�b�r
7^���|�+_��n}�m�h�������Nu,���!�=��]�a������lf�D�\:��6���OeHx���={���g��>�����݅�;�����pg���V���n�
ȕ�W�]��x*P�P`��<��g>�Y'�b�_��BO5U{C�!�̙�1�&('x:<g�X�����wZaxpD�FM�g��5r\|膁渖ok����"(�����4u1?Xo�������q쑱Q_�:?���D��A��uk�z�0�����gW@w���p�T�)�߅bֱ������ׂY�z�:[�bC�#I���Q	�:��kϟCDn��0��a�Řbm.J+�e�8��m���{���ҿ��;��!U�q�5��u7��T3�^z�S~�C��1�J)M 9��_잣�O/˟��Y*XU͸�ᡟ�:IbU�����^5j�.X�<:�z���C��׾����v���C��!��WJ��>��hr�0<(�U~�'^�^	���C_�<X)�ël��~��{�}v8,".��N�F���cq�g��i� Z�<6@���kEB��B�@���?��@3 m3��=z�K^����@�c5!�9��P(T,u���a� ��)�a�y9���պPMVd53W�)�!_�� �Ie�o���qm(+<<8͕ J��v���p��;�A^m���C`p?FǆGFI��������X�Pf����7����\8�ڱm�Si0w�k��͚R��<�_o)*��d�cࣣ+m3m��(�f���n,�,,��0$`�Ϭ���W�Q$cH-�'���>�g�� 2����e�U�ׯ%<�o�sή��
��w%�F���O}�� .��i��o{5��?���v���7����/�3X�q��:��YK��_����Um�u�o�� �&�R�88¦:v�MN�� k��M.��x����8�#*`�QYs����y
Xt�z)��u����EpO���-�u� XA?p��V0���52~���;|�#��H�r���2E��X�m'����~�y�#>���ѹO|���� ����[�l��,�Ga �x&��s%���h��q�5kW9$ǳ�y�]~�����\�q|^Ûcsc��9#����(����!���k�E����-QT\J��̱yM� mjR�|)�n��5ǽC�n���Y?NW�.��Șٱj��{	�V����q7��m��I�J��P ���{�)T9P��s^�a�7rl�F
=��]�z��q�����=��ɣ��r1��k�s�3M/���b�䄑X���������.��a��+��w�;�����/���gݶekx�-k�j�#��7^ikVӏv�ff��=�`eWmo��4� �og��+M==y�~���E�B~N�K��K�sW��)q�b.�^����j�����>�KG<b1/}��Kv1�VӨ)����'%KU�(�#�Dt&FL�����-�"����/ӿ��Ω"�p���J�yFT�JC4'������;Ne2BQ�Xxfs��~L�;׆���t���N�^���nܜ�&�0�3�=2=x�(
Un�lX�^tA @����}�QkD�+�{3J�/�>;���ZA` ,/<��銻}��6;q�S�[(D"8h���aO��ۥ#v�nŘ�O])��)���;��k�u�4g�A�¡ D��*>�z���Ԥ=��=�rŰ������#���v�G�R*ة'��ذ�B��}op^���z�g� �z�_��Rtv���XN��� �N�,����a�@fV�F.�"��v=h�a���dP#���Q�?��?�M�Pb! U ���Xo��|_��d!(K�x�Ҋ�Ƭ�*0�6�њ���ɰ ໯�p�.gt+,��l�B�yh������]X� e��������X�,�f�����P�\;K� �5&x*J�󲱸'p�K�=���~,0��g~�g\� ��g��fR������[�ͥ�s��=�v��
�d�_6=�k��g�ry���kF�?���v%����'̕��@�̵���kc.bC�U3z��2a]�X�W�s�p>�g��1pϸ/jCyn�QH	tm1�?)�<�X�_u�W ��=yb�V��|��6�L��I�pK=���l,�6/eee1�Y�@|�4s����«{��{l��Ƿ:�g�E�p����S���0�B,���W�<��̉���?�y��IY���(��̔oڑQ6����A*�U,Kl�)��iz�f#�T�u
f~����R��y�b{!��c���9;tp���}oX��66^��k���E��@YZX�۷�#C����+A܁�@F��E���k\/��DM̱���5���N"�k������:΋@�;Vp6��c']�#�Ԝ��،��^����.3s^�zE313�XPףt\^G�)~�@�o�r繂���|��Ԁ럘��������Vf���G�P&x��ȍ�qn�w��^
־�1��	؇�T�8��i�FA�5.͖w�b�;~Ć�ﱡ�UaM�[��{��k�#���S�����
��������a�������7����z`Ȩ��Ӛ���ke�(z�d��"��"�@��b,qxd��Z�"W,O�"���)��>7��l�]]Z'���Ց�)~=��K�r��[��7l��%�V��p[�l\�����?�������\y>wki^���e�?l�sAIET�3g	��E�(�"��ur�[͠h,X����u�0����H�s���j�
V��/pKA�2�
e���~b#x�pB8��`��^�ʯ�?~��杺���[�¬1W�k���.�q������#�jժ�֨ovܡAM�/Ͻ�9. 9��ب7�n4��ޭϸ�ߓ"`�dg���}��ܺ���+"$�7�.Jx��5���O~}ܓ���%�l|�F�m����k,���~�w�r|��Wlz�7���;��B���r�����(��[�9d�<Pd���/�y=�Y�v����� EI\��0/�~AJ[M���<U��0�RC��& Ȱ�qTӡX�֧��i���TťF�!���� �뾐d�p�[����xk{k�T�e��1[��v\r��׃< #���S1hɕ��q�Q�����[�?��'��\د����ۯ�����ҋ/� �����)��JT�%�@���Q�t#�X��t-�W�@3�ylx$�g�T�K���R�y���j�W�!K;���vX��9�k�{�iG�����w�k��9�U5�E����ի^�P�0ؼd!�����j+&�Q!m^64�D���>;z����e�*��$T�˖�B����Y�g(�
�m{��^
 �}bO���0	N ��և4����pN��9�Q�/֋Z�?�wP��,&yBx�2�a�s��fD�'�+X��u|�s����C9��zZ���1����J�L�5悧!aԣ4���f~��c)5��B������.�E2o5@W<F���Ҋ�MxWR�D�K��X��� ,]JR���v��z���PŸ���R�.='N�f@�3�^��sL\����(���8y�{�T��'�Z�S��k�(_������B��~Ϟ=�'�'��׼�[���-o�,Ω&���W=ﱆQԫ׭��bSӳN�7^̮ەV���ȕ�e���Q8ݵ�Ϡ�Wp��b�7��W<88����_���pݵޡ�۞���C�e0n���uހ�߰2<Ԫ�;p̨�A����K��y���wz0\�\v�BXW]s�o~`m�٬� kyfz������f��m��a;9=���iD��r\� y�r!�+�y��~C}dU��o>?���`�"�����`��]�U5C�H�_�zsU>#��&���yO�T`�X��6���P�����>|�M�5�y��F癨Z�g�޳�_躽7l�M�1���|�P��96�������ؐȫ�[V����^�PR�Zi�8	"Yв��B�@SN��	�*ӊg�ȩ��e��U�:w���ɭ~>j�����c����W�Y�4΁�H�H%& v
���DY�z���H�W�4��eu7s��\�X뭬��@'�?��'&��|���.�](؀��2��=i�&gmhxܠsvt!�Y���7���}�+�؁�/��灂�"Y\��H���"�L�.9�Ë}߽��ϼ���Y�x�6����AV��]87���[��E���s��n8>�?b�T{F�Ӽ��O+6�!��bx������+e�ґ�>�屑!۾m��_����:x�<�a����CA��=�U���BV�������.�!m��K/w�W����&vh&\#�3B�F�@{�	��`8/�
�C	�0�xE;Q����3�u)F�2�\�36PP0�	e�<H��~��x<���o|�=���Z�(pu��N �{� g(�����q��|�����/��9��F�=�<o�d�[�� 歴����=���=�뮻|=)�V7K�˛J!��}Rn����LxJI�8��RPEw
󤰍��������+�,a��+���-��!�+� �=X{����_�����a��iZ,�g�'�{�}�^����~�����R%�ͺ-�o���@x���<P��Y�����u�:�sb �Y�x��o��M�k��|l�~�k����4�A�tl�m�y�%���M604hS�s����B����g��_  �f��j���ȋ�O|���[���m�~�w�yd�^۵�A����+H���˞f�_y�]|�����qc�k��h��_�W��y�L��E/z���%
�C8h#�z�ڂ�ynz�>��OZs��!-��1����5@�<������`��]R��+��źP���z�k_���?����� <�������T4 
�J�K"P�%������Cyb�*�&�0L���tL�/�D����gȖa�!Xو(���o��m����i��{,8Rq�\?��?�0X.�h2}ڲ�Q"�x���.8���T�F�=YK(���7��9���7�1���^ )��e��%lH��f@�Eֵ�q�P��iuu<y6�w�
l�C�N���dm��.VZg2���{ �y-���?6e*���ݳ��{����A91��-/_�6+mbr�ceP����;mF�����'�vvO)Q�C��d�Gq���+5`X7�x}�C�֭�b���>��]-W|Τ��_�=�����z�&��a����g��q�q��~�
ݚ o?˹F�>��Ϻ۲��`��ƛnJ�{��~��`�+׬���.�e�"��E� ���ᘈ�������rx��a��Y�A!�$��<��wx�w�=_����`��:�!�(�u>zl6���rh!�Se/n��>�-/�1/��Qn=�M��MДkG���6���Kγ 12�E�	�b3pl�G�V$���*����̅{I�%n/
��3��=�H���B/�����;��fnT�FOf��/ރ�Ұ�����`����VQYH̓�^k�B����O��	b�S��Ҩ�F��'� ������[ǂ�u,>�='�h�S���1�*W	qF��W,@�[�B0����Q�<C�-o�����[���ӟc��1[�r؊����ʞ�I�;�=�5�6���yn��K�o�} yld��R*�'�w�?\�!��M�X^ׅ����FQ�$���Xx��֯�U�/��n��[w��?u��2��o��6m���0�w���ѻ?����+�Y/��ֻ�;�T1p��`�~d��ٟ��^��Av���k�k���HŬ�:��X�ln�VA$
�)��`RV�\������tK�E��������w(
B����Y�Oz��T�f.;,�/��S�V_�e1  ��IDAT�9�N[ذ�������
��=��3�&�
��,|\�T����@�\#�8��1Ҥl�(�
!���Ȇ�ް�8BOE���Gys��e�f�R�����h�3�g��E�rI1rY�\�,e:�����~l��!�Y#|��B��s=��ǣ��Ul�$DdK(J Kp��K(+� ����
�+���4{DB\i��e����|����$#�y�K橸�2�4o�)-EvU���n�Ev��WS�y��V���gf���[��+lj���1�|h�X��O*���tO=#�򛜎�is�>g�췗������~��z�Z^EVpr�{�����^��^�5<�<X�+l�E�mnfֳ�FG��.�+~�#=�ȁJ����9w�8v{��O����N�� C@��Y��@,�w������n��6�,V�ɐi�,��Y��>v�G\`i��0��@����q���Y��=�x�;��X��%J�%1#E5(�JǙ;K���
E�}
��_��]gb�D��oȃA�2#�	sF���#\�����pl�9� �V�ŀ�&�{bGDx��;���?`"e�7/�����: ��6B�\z} JE�[�����r~�q)���
��X��^��;�c.̕�t���qߠd�C�,��3PSp���|��ZB9W�U�Pe�p-|�����P�fjy���R8U��"0�#�B� ��#��*��uy|(��� ���y���k�xf\� ��?�A���c����8Ć���}�T����U�"��{h�f�Vۋ�ʵj�������E��@V�u(F���5�������]D�X�y�S�[����g]��-��]���62dM0̠�����=�v��G?l����3�ckiI����6��ހ0�&�ed�<�QK����}&XjP ಣP�G�G�Gz8,��f'���k�"E� ��q6�d� (X<��ۿ���i^�R4�u]YMMUm��	+���κ���wߧ��r�c}���c�C�{���@8^x�_��}�V�QH�D��9�"�6 �S6,��������TF�
������
G�1�!����B �>�dc"�`׽��r.�P%�|�7�e����>��7��
�p�@ �!�U�P�?�˵s������b`�PM0W��'k=%����d�=��FW�X�y��,U/�kn��V��ز ���Ǽ喙0�geYO���{)���=��e8ʑs��Pp
��.�4뽖Ѧ��R������_p��l����ɪ����2͍���)��[#��s��ǗŶ�@��Ś�B�}S0&/��J�X�������͠+ŮD�r��q�����,�L7���k����` pe�{�.?PQ�9�5 ^Љ�]j���
��?�!�{��͌�˩�x��	�]�ͷ4,��dq��45�ZeC�`�������/����O��
,�3�����Mn�⡽�>,�^�V+�>��.w���-.��5d5���E�@pE���:x�+_��닻�)k��]@����`T������T����l~��jV̣��:J���	kW�+c�%��W��7�r�����ͼ��:O5D�U�&�e{`щ���'�'�G��֑��T�(�+����\���&����J�w�f�Q���hrr�_S�XP�j�Ny�"!�'�|��"x]�(3k���W�*2���L��u�
��B��_R؉������kG	����5����J��u�&[�vC�C���F�f��2Z�ڡ����=�p�IH�0եp�����T�Ǌ��=���S�>�;*ume�Vx
"����no̿�]�'�]�5�e��Q24�7>ZT��B:5�� �X>���M�<��M�Wit���k��`�u�b�F�����Nc�n����pz:����H�Q�
T
���B~��2L�`����� ,��?P,@-Ef�Nf�7i����g�0r�<�ShcJ��hKA;s�ֲ�����"!��+y��z������*|�^H8����dR�^�J�F���q}�#c�-%����*^W� �3�,87�e��=��o{�E2�����`�c�
�K��p������\熍�eW\�ﱽ��t���=�����u�����f)�<�/$,��"�U��i��vs>�薧}�+
�#�?I���_z�Vw�����g�#>\��Aq�U��ǟW�]�٨��+k�_?���Ŝ��=�=8������xj���6gJ�Y/����q�t�eeҼ��n{�MۚO�K����nXWX���z˒����K�Y
��z&+����)g�B��Uv`��� )�>�8�AX0X&���gr\�,P M�N,<�U���lp,HÁ8��9��8J`#ă/���p��b�*$��=T�
�HlŋUJ��x��z���,�� ��9�I<�(���x�9�+׎@d���/!�g�G���cP2 �Rذ�|�����ٟn���z3��7� W�UB!�V��WU��2uXlz�9�Ph����
v#��\|����s.����꠆ף �<�����j�9ǥ�u%��5_���+��ݏů�n�#��9�ei�Sa�<��=�z�Iߠ{h4;q��b@5镲 ��t���)���?�'�5�<P*ts�گ��BLKu�"�X��sc������_�a�g�-�j>�E̕@K$K����<�����))��=<,R9��~�^���yF�K��#�û�M-gF�5�"��W���^2��,�Y�W�&��{�U׸ %�K�
��I�;���{�\���Gq�7	���0J�+��Pmx����;��L}�
����h��LP4�B���rl�N)�B��CJ�� ��9�
����5��X�j�5�f�w������,���

�`�ū̚�j5� ����x���� +J���2�!��0�W������7����1�N!�̑�@�F�P�iL(BYJ�-o.b�B�F%��'���y�*�z�b&��B���S
�̯����ql���(ԭ�l)�<���B���VF���4+�LZh���U���`�n�/�p��m��gPP����c�I9) �,��^@�s�e�� �2x�E�����F����������p.\�au<_�=���l�ѱ�3x�:E6E�S������M�/]kl�"��d��ĺEp��!���۵k����w |�4W�늴J,o�K�t	*	8��c����y+�4B����_A��H�D��u��7��F�� w�X�j��2R�s�-�5s�(3���ÛA90v*��!�D_�y�����+~e�(@�5�I��$P|�&�7����hE�Y*�|xA�?���\��E��d��� �h�����Y����\}��2���,.%υg�ץ���'��f��ĜQ�<_M
�i��"�no/6�]=����Bs�p�C��U[�:�̍���9O���Պ�n�� �<G}L����5������T�d���h:��E���0�b�9Z���?�������9��3Y8< ϭ.ƻ�ng<&����Sˀ�|`2D�'#b3w��  �c�%�=�J�;q���}Ȏ���
V!V6OS��-�O'��S�TQ*X �4�a����Z�H�!@����4]EFlz�� .}>�1�TʒM�<��s?e2�F�qQ8X�X� U_^��\�x�;�ax��L
#�J-�\��5�=�X�y`=��B��� �a>QAY�YLɬ vz�h�z�:Jc�+u%���c�O��&��5 'I!��<A�xR�>���m�>�_1Y�xO�o�פ�Vz��I�H��!�J=���N^���w~�b�b[�Jl{X�1��	*����.�r�_#�V#��Y+-��n�'U���Ih����x@�qnJՍ��R��]�օ�g":����3�.�g���������6`NY�-��}ou������W�7��).o_�5�$ L���m��p
k����c�lr☍��j�#�2�}��+͔�gyZ�!��<�����o�'m���%s�_�`�>��Kإ�����"l��:�G>x@-�!�!�KU���e��"�
���!��+���%��2��`05������ �X����=�n]*fJy��kd�xR^�zRПav����L��!��)K���K��Q��k(t�T����������ͣ�"�w���3n�նl�(�����~�a]�ךd.ɂ-'�l)*��g��]����������9���٨ (ҀX�N��)���nVx�S;Ik�">ǉ��{[��	߲��4��h�W$ռ�Q�h�~�w�x�2:a^�v�;�6�E��_7�s�ȫ7��r2��S4[u��|�U�q����NA�,�>���i��$�ѣlwb�03�T��5����A,���p^]y�l"��XlY}���V�v��c��J){Eo!,�f�b���=��٘�e���@�|A#�a�#���������6� �p=�{ѵ�]V
!&]τ�c}�#OP% FL= ��e ����Е)�Fձh��|�ǀ@�~S? U��ൠ����|AF���I� �@m�><M���L�Ac��&hG�>ץ�]�,�@x��s��f�(0�BF��f)\���0�fI	��N��Z�����ܴ�����~�ɩS.\f��5W*�zZ\�
p]k��n��sn���W��� H=)6�Ou�4%��$:����t�3���m;?W̕+�
��O���^~���-W�P%�ً��'B
u����=/�?35�ߋf���������-��{����F*��-pE�9wP&���t�)���9�X���x}��۹<
���k9�D������4#L.ndi�ܞ�8�F�"��z-���*���)>����^B?��+=u=a=zd"X�E��� h�5�A67\�z��Y(s��7�6�(��SgScR��,0	8��.X��M������0{捀U����P�g�����d���je� ���̊���s`�@7���~���>�<��96��<,w	@��T�)m����A�)�ϛ���R�����86�'�+�WZ�80��ԪR9�R�R��$,w\�.*�ytM�:��w���o�-�̇�������yC�c)���3�"D�\�=�}��
�����kIXCs����y�
r�6@���	�[z�L��,jf6x/��%��9/جt�г٘�}�w�Z����>׾��1sϫ���(dJv�R��f����7F�e�s��'O�c���#p���-,h��N	�c��Z�:�?����oΝ��;W����nӘ��3\���2F�%�.h��\�^5k�*?l�Us>t����e' א�'�[A1Ǣ�D��t�?�͖��x��a�
�xF�\*����U6[��M����d����[x��s��s!��p�4��5��'Rl�G*]/~�	�� �W.�R�<�e�I��}��bl�����	���X��A�my���,�f��EX����+�y�0�����S�B�_P����B']_��jϿ����#s/4[+��S�H�&��p&q��<#�%�;�����{�>	x���(���Δ���bAZ��պ��y;�W�$u��IኧI�N�������&[����{eͶ���q���M���N�\��{-(�L�1�b�i�펧���?<<j/{ɋ=A ��b^�������9J��^�g+�@c@"W)Ÿ��̔{Jp�7W� �9o�ĺ���q��Ɏ�_��������j�@�}����y�V�:d�@�w���BD
,|Y<
���O�X�T����,#B�-�������Q;z���;�E,�V3α)�FƖ�l�aC���A��#�U��֏Z��+g�4�X�??�@6�|^�b?�-A.�T�\�Y��LBL�.���\��#!�znj|�"2e�nR�+��\%����ϊHB_�A�H��o	���ы����(��*�!~bg�Nn�ׯ3:����J��/IC�&	e�-`.>����{)/����o�)����Z�B�����C«�d6q^���`z&�D�.�
G�NJM�a^��V�z�s���a��lnf�s����䐞��[6�Үw>���g�
8Oɔ��o�s��L��=�g؋^�b{�[���.�w���5���ZԞQЛ�B�əY?���k���$��Q��r�a�}�p��Y�7�Yz���P��*@���ew�U�r�j�`�\*n��_�����S�G��6��Y��cA�o	Yy(8����`�B�~�{�ч�e0����Y�B��g��{��y�a���K���w=#������x��k .Y^�Aۮs�p�'ON���H�јuET(�l�ju �{�s�*�X���l����`���BX,�
�!��Ț!HŻ�e0J����}�;((6��Ș����ȣG�g��M��S��>�h���e������ �v>����j�=�� �)z�(ޗ!�w9���k���0T`W0�`��������e M��DU8���9��;#��s��/���ۻ�ֆ�T��D�c�i�P�C��p��GF�TfAn����3J���V��@,�����n���Ea���Zv�����M�=�r������}ͮw�r��(��|o�˷9��1Q�P�P�� /�����(C��L�FO(���O:/��7���8
��# �Y�G���|���E1{	:���3��H�8G{�v�0$(����Lx#t�կr��a�V9��Lh�Ć��sa��'�&lU֭�>YK��L)�rs, �@�.)�i�2��j����@�.��V�;l��I���]1��`�ݒ�x��>+@�L���K.��5(���ov�"�2H�)��9�k+%S|/d�|�w=��X7��ʓ�(�����$%��$0xj��UK��%?�E�%@�(YJl.��$��&'<o�2!���,|^�:���%e �;�Y�E��?�"��^�qI]�>�*��<H�Խ��|��� �h,t�di�����}�(��	]�&�&����1��{��E�0_�����U����K+Wr1���mr_�kN3�� �'*ϰV�\�$�/������^h��2������9gqu�C���(���LLĊhkG�\����K�-˖۝/{�C��aR��c]��e[�f��ر�>����������A�]��ȓg���7�ǣ�x��٫^���za�fc�EK~ �~tt�Ɨ��-�0�*h)��1ɒa����E"�EJ0T<X�l`�}ua�9=.���W�,�bݩ��S,�4����\}*K�+�5C;�6��aS�ؘ󕅧�m��s��J[��2�2��AKZ%�A��M�~�(ā��E`Rp%:,Yb(A,"�K�'J!M@�cq.�T�у���TL�� �Q�(-�[j.�0`ŒWz(���Qr=	�r�Xn;�����,f��=�؍�B1�bD0���W�<�j�@��z�����
e�\"�	�4՘!�ε��P�j�.��X�֋��GZ4���j�Y����/��/�ڱ����x���;�d��������f��1���Pg��;'�,�P
JmOi6��4��i�}�I�+*��h�N۝�M5:��S�s}���� 2SN�Y�O�Ӏ��oϞ��>f�)���W����ړ�K�-�hX�ϸ�&�pi�hjjjL*/,c��j��9�U�8���)oϪ��Of���!�E�f�*�>Y�j�����{Ͻ���v�����Y	s%<��o����&o�c�E�1�"����&��g�gsܛ�A
".$.6��Rz�F��U���r��E]O#]�|u��5fO:��C>�*yJ�Sp׶P�Խ��W!��(�兒�|���UW�k���9#�j,N&V1����w�6%��M"J�h=E�%��EѢ8�.
��x��PЏ���pN	p6$B%�����h��$� ��s�������>���{'��MLsn��(R>U��w�f��1�dF�b�z?�M��:@��ޑ�z���2\R�����Q TEE��S�Y���KR�1��3KV�iv�Y�C�K��7J�NuY�:��KMg0�����H�����'ҘA�{�&&�����%S��$��
{�ہ�o���.'W�+|��J���
t�{�A��zXC����x���opo�����"��P��g�S�K���v��kS����#�/���o�kxN9Lz�u�������{1zX���G2���n��}��;ۇ����A�_v��v��O3x�[A�۳���_m��a۸�r�T���%���gϼ�v��W��@`�R8��J��(��Y lr�����l����-�4�s��-($kl��m�z�f��>n���¼���:O��w=��sY������a(���a�b�"���" �0X�@���{jW�k�@�3 -�{�E� ĺ>�7�e���`�J�?c�ca�T�~���Y���&eǨ��������� #��|�NA+\�j�9�h�sǺOy]t�P�<s ��84\B^V"
����?��� ���	�WN����ZZ���k�Z�>(k��9?���Ȩ��f1��S�ǳz��_�`���ՙN1
]�e/��4;Ią�����1�`���}���U[j��>Z���(���6ۚ���_a����C#nu:��V�I�����E��� ��w|��W�Ws
�=q��N[�ض��v�׾���
�t]�+"�i�БÏ����{�9w|��_����M7�b��~�ב`�T������/�����ٺ����M=����o�@�����8h�.wpjj�N��6�χ>�A�x�� A��sYQ�Q����	k���X�i%c�٢�z���b� ��Ҵ�e�e�k�7��2�x��0��sb���u��ӿ���֪Rf����Y����9?�!�U�L,{�9���_��s�4V5�� �ʔ��ō%����gs!D(�����a�X��<���]'X����y!��c�i����!��(&��uE�9�r�y�¶96�F��>����R��+HY7�(�aH�������7bJ��!�eaQ2�0Pe�}�e��:���a�k6����&\��;����2���dw���\�,y"��bAٙ�Ӫ�Փ^
���\;�|ݰ��s-��+�A��|{��[-��kT�chx�"kUƑ�Rd݋J�xz~$LM�8a�����o���p)��:�@��������W�x�����pҳ�%���i�w#�Y����T��˯��Ղ=���v�U��E�օM��Iϝ7?��u}:��e;����?�^���������\$d��ԉ��#�x�q�Aq�����¢��y�>z$w����}��[KV*EXyzZ1rxƍ���Ѕ3������rJGeQSEK�
x��d�ј�t��",��jD@#0�,BP]�Ԏ+�{�o6B��`�# �Q	�b)��S?�S���"WC!a�� Q��&���?ޘ�����X|�g̃2�k!��5���� ���>q� "`%�2c�\�ϱ��|��5A#d�p���)��Y��SS��+�eq�1�Tx:�JMv7/��%��En��o��1x�z�|�9I!�90g>#8�g�{|�S��g\����B���9e�Ⱥ��`<��G!YۋX=S�G���Z�زѱX���oY�V��`q#�wQ�ԝa���>��v������*������/��/�JC�!�x�x��`կ�fk¦�&���.yOP���<�^��o���*a��\����zљX���^����?4<�س;�s��:d�`={�CC1`Y���Z)z��MDe=��c�n8�?�s?�.?��B���~��XlJӫs:�?��n����O�KZ�d����U31y���3J�
�T%��$��9"�����H&����c(e���0 ���AEW|Ndp|����P 
�i��5`�r<��#�M-�2��=W�.�����w�����( )60J���#^�Uv�@H�(M�8�l�(�h="�Sȱz�S�[�4z�tXk�����=I�r/�)�9�p�0#J� �o��o��������yQ<�Ng��k����_��1GY�o{����\?�Hyf��{�r�5xq�K0���<	�`�s���y�y�]�(1=9�$
��cC�A@�O�G�@Φ�A9�xm@ ����܌�{NOO���
+Vm��q�dDF1#O�n+#v�gdU�&����1o���|��Wݐ�6�}�q�;d{v�
��B��jՠ���(�:k����{����r�3=^�^�:�}�b8Od����zc�1�]8��kqC� ��ix�O'X+v<ȄU_�2UySS'�����0p<��(����TH� p�����1�(-.�⧥�5�_D@O���ܢ'C���R�Y<cˣjV�> �P�i��;q���o橬���4�F�^}��2E8���%�l�3���6m�����íJQ-fq��`�����)}!��CmJa����b��+���ڎg�}q�W��ann&ǳ!��ξ[�J�;,L�x����q�V$�	]�=�ɿ�ï���9��������y�A���=�;�U�R�+k5-��9���y"��b�f�i�0w<�>���|�Z��
k��Z�
n�[����0��۰�yF#c'�@��ŋ뱩{��J 7�2���pY���`y _w�e����ed)u��g4X��@�4O�si��SB��g��r���}7<����~-v��n��
�X�[���!k7c~8<�Q`�S6��i�k�"��[��X�0KY�(�#p:0oa����h�BL@D��|���\�N��"���`���	�F��h6�R��4��[:��7�*V��)+9�#��kVPQx����̊"A
D�CA��V�Q�@�nZѫ�p\�V�'������[]��-*�Z̬�
`���ôЌ����֐�"�b)l^�󋋲Ty�Z~�P�������R�(�9?����MF��5�y��&���-�����P�����Z�x)�/J઒5-@C��$kIy���=�	����ow8�,1�jyF2���b(Z��w�M�ܵ���}�㠪�j�Ra��,8�?���G�v�X��Gl��N��iv3�:ˈ��N砤����l6x.@�p�?Yh��T��5�����+�jPp혵�=�v�Ѻ��1�Í��P��r�Ki�)�G/��y��!��y���d����A���j<�bL�D�V��)
5���c�P�	$�xpP
��	:;�!qq	b��>��M�⽲p�������c;�՜
�aN���i`�x;�zv���]xͲ&�=�(�S��`u;'��~	�Џ,e�H��yT ���:�\|5�Q��
�Dɠ@eJ��V�J���_/�%��*���)%�YB[��g�yu:?�PE����=�L�e��6���C�{!������ҌyaĚ�b�I����Q�T=�Y�7��ҕE�̓��	?��c����x�<��=R��A��ʘ�:ԁ}����K���"����}V��<�F�!�9� ��e��8Vu����X��O���m�v�� �n��w�\�Gcü���±�v���/5�W}�x��5���� ���(v+�2��ky�������v�8����������)���[zo�¿'m�,@��b��kæ>f�\|�ՃU276aa�jU�
�j��D����h�pW5��R�X,l򾱪�_���zVi�X��nq��M!���`��)=�}��F9�@m�f&OXi .��/D��Sh��螮�E��@#���|QG�k�*S�*�,��զ�q*�9����ɛ,e��m��;�D������"v���)��M+��{A*���'˞���NQ�oR����b���GE��x_�E�:X/BP�|GN�R'SG�S�'�R�j1NDy��!6J֯��xMp�FZI���EV����hR7�Eʇ���}5�)��ސ��Q
�7<%��p]��ĝ�_ۧ[���Y��X��	����7u��k)V���O>Go\�)�궜W+�Y���;_~��Q�"xU2��A�P��z����X�p�I�8yȦf��h<{otl�O�ѵ�[���=��9���h ���@����R���/��pn�G�n���%��+�28d;.}��~t��{�q�/�ff	tl,l�Ma��p�[�v�?��Nz[F���f�0�ʀß�?15i>������ٙ\�a�PQ.4��m"��o|�]WT�2�,�Y�p.Ulr�aA&��ȐMM#`��מ�b�i�}1�SV�E�()V'㪱{,,Zܩ[.8F�E��+�@l��(�=J3��L��������"}F�KiR�Bp�vJ��ІO��H	�t^��8H�C
�A�Y-R0e����|�@�E��\1�w�	
c�W�R���~��`������`�y���2�39硃G쑇w�.���*e{�?~�cSk���H�կD�Gw���"{��̯����mϣ��z���|�n?)��������>�1���
�5V������e�:�������O�/,:�w@>��OL7��)�mv�m��T-�{�1��I;r��a����t�^�5��K-���$7zPTp���C�R经��e�����=�����<[�9���m�}K_�re��d�uY�-7�Ɩ�&���m������&�����1[j�K9��˟�\$C�v�؃>ܫ�A��-��ԜW��߻/X���۾u�W���;qrʭ%pU Ua]���X�XTy�)���"J3:XLT�����qZi�܂�:2��`�dn}7X1mk461�p� ()�V\�7����J����к�BM��x�J�����R:x���/O3�FA��6+E(+���N{3��oY��W^�g_��)�df���*�:��C�Ǩb7e�1��
 ާr�c��CV��`-f<[ɕg�6�
�Յ���k��u?~�F�3�{ ���Η���V��}�/�ۺ�B�Fl��v�ȉȔ�U�
B\�v���b�����dT�Ѷz�ӥ�LƐ|����>�����F�e��I����^���UNi;kW<�Z_fG�ǵ�v���~�F���9�m�sX4XV�?�a����A��X_4W%��q�I{##hn&�2�����߽�A�������
��@���:	�em,�����^�:aِ���??��C^��7�´]tA��k�� �`�S�@l	�
�C��7��qA���H���(�B�ě���<(�{��R��|d8(� ؏��a���SRb>Jc�����?��n��\8�(�J�U,E����<�y�.���LA�³�÷�>���r*���&�0��۶^l/���Ju�9���q!��Zf#m�?�On�(���`�K�*V��T����v�R�g|��mlt�6l����똚8�{��ͷ\���ꫮ���"�C�'���͹3b�\j��¿k}�8*�&����{��?������k~��ʾ�m��w\7`��G����#I�t�����
���l��A,86A$gY,-|DiZ.k�J��yN�<<6��I���U���������d=kA	�J��XP�Ƿn��XZ�J��uKД�F ��k��De�G, /��18<�4&R��_�k��)�f1l��L 7͒b�Aq�7���]r��8��ķ����e�(��Q�U��K�}%�Pu 1!Ȩ�`�/:<K/��m[!^�f$�9d�ʒ�1��_���;�3]��& �Eߨ��}�?�Ǐ����g��Ipu)��`OWka�+3G�nt��k��=����l�5�7��-+�ݬ{.�<>OL��ۯ�{������Ïtء����=g;y������I�G�9�!;v�����ĭ(.鞠/��%C�u�����ұJ6��4��[�5�UF*x+/X�,�i��a(ȉ%��R
�-����*2�_�5kW�f&X)��
��9�aSԃ��n�*�����Tc7�蚗=��������4&� �A�PP��5(jkՙ`m�D��&댵�\�X�.��F��J�e}��N�=�¿�c���0K$�TZ#�t�K�{Zl��S\p^uv����d�n5�Q�r�@��g�'K�Y�1̼�pMk���.��r�`���Vm�ӵe�c����50�}�@'=/�����S��?�u.1>��G��j��P�4sQ��I��f� >���ڱ#��Ѓ��[c��68�6"�Yg������{����X���=����Y/��^��0{��ĉS���7�Nǃٺu�kjR�H�"O��*�͡^���ȌtNh�y��M#r~�|Xboy�[���H�� �U��1���
k��M�)<�x|��a�u��bFbN I��,�X�|~|���.@�X���0������ e@!$ș'��
�2߅v +{.��9>� ���M9\T_����W�@V�����C���J�5-�c@l((�c�߷϶���^�ĩ���^��AI�'�
H12*��^ĐY�V�����=�����͆�K�[τx=x�����F�!�c�p�����s��/X�6OTP]C��J�#����z��:�@���l٘�L����p�=�e���C�r�������l'�~E^1x��ȐkV�W�?��a�~���9�m�k9g?��MF&@ڶN�����]'+@�N,!�m���)�,k��+ћ8�ųe�6�eu(��G���7i����N�5�_*���`�Ȳmx����J/L�۰�y~�|e�Ɉm�u�Ќ�M��^N��6��5mө5�{� A^�q�7�<^���C�����\����<&�@��7�f� ��@)��0g�S�
���O�U��b���=�sq�*�3{�{1���"ݼ���k�>lr[��0s�T����g�Ůt1[�*�B�p�{�3���&v"��稩�~p���磔g�~�����>�E�r0�����h�2yj��aϊ|p`8��`?�8<��
�sS���Mr�dYɺa�@[1�փ���j���E�r�������1��Qx��%� iǔ�*��HpG�l��6���w�c{}�S0�cp�K�c;�J&L:9���4����k��a��!V�z�:�8���EN�ų�b��HM��5�����Kҁ��-9�T���lԱ����w��e�h�^_�җz���80�x�"���5��]�g
Ͳ�T�+Д���u�*�4�3����C���H�lWk��y�[�nS��P��b�K��xz�Vu��<n���*�p��u���T:��xN�� �r�ʼ�T���^�y�{�{�.�(��^�w�N�)^)|�Yz ���P'��[���%#�F�sb&-�/fe�N�fy�_�b(o�EΆ�J�5p~�a��}U*8'�PV���uc.|�+5��+�A[�b�M�<n3��
�����T��F����ٯ���K�D8 �`�KR����T ȿE�&����`����վ��3��,��CL@5(	������{�;�5���u�`�°��\`�:7�Tf�F��\�I�~+�o��H��b�9{�A�_�i��[���!�2�T�����#�S/GM
�R�c���m�2h'��AM�u�����}�7�tP��*�3��ꭺ����n�"M&sJɤ���(�L�������}V�>ޅ��� o��B�4�Rʷ��B�"��&�%�M��w�����:�H���q&&��Z
Mͳ�x���݂c��^��ѷ3�g�V�^^�Ƿr�/Y���
_�W�g��r��_�,�aQD �U�+�Y���`}i
�x�u���f�ȏ��.<Y2�87q+���y>G�&s��L�}Z����������x-�̤>~�K�8���ڧ��e���]�:Ԥ�R(+A��	�P
���v�N�H!�L��lN�c�O��{:7= D�!�������E�O���7��_8�D����WK6O��0����yZ}��7��]b8S��X@,l�XNlB�(cH�/�>�g�8�ڝ�X���d��˙k�ͨ4��Ջ�Ƿ|�x1��@(L��Z-�9.�X΂!����W��pf	
�S,��ǎ�m����>���ń��k�����W�5}z�}�Mp��H��~��6^A ��@U��b�]�X��&p>C!��Q'/)��A,�Ua�|�T�(/��N%bX7p;�X��r�t��WD*Z�V��ͨ�ݓ�#6T�g�gڍ�^,+R�g�z��ݷ�H���߽UZּ%�P����t�z�_xB����|"i�����v��t*	_̕�,
����S�8��#v�P,D#�'6���I2O<�y
�,��<��m=�U#��ֿX31��h� B@�����x"|�|��e�� %��Y�+_��(��k�@���Y�{<a��+6!��6�|��VsQ@$�b�s.���!
׈��us}�n�����Ҍs��-K;3��GOZ������И՛���NKy�q_f��ќ��p$U���PBJWr�C��!�o��}��3K|���z�U\Z����Xe����HcbStr��f@���g����]�}�6[�SCT�5��>u�U1����6�)n�~�Db=G�f����0����!�	��u�]��?��?��yV[f��8�)�|:r���g�������:��Fŋ�,9��S`]#�	�-N@��MQbc哵�<$������ �`�������z!c;B�Nk{���hp�?�����;.��1}����=�R�
̺1�윘f��+���b�ǐ�#��Wa1͢��su��q?g����ȫi{č�ajh�*�Gd`��Pڨ�r^�q�[/\3X�O�ɩ��lLY�B5�y&C'�T�f�K����dXv���v�����������3��e�,TQ!���:R� �bS*R���pLΑz��-b7Q���[�kJ{�w�J��G����`G��Ҥŭ��BOEe =~�u��.�0�V'B�@si6;�6u����e60X�L��R����S��~�=��RA�������k�57bY�w�l�'����	�?װ���,��h����قֆ]�*%��!KFCʡ�i�����ڀ9�s�C�Ϯ/^���<�Y]7?f�0�Ώo�L	Q`���N����4ax|�C#ܜ����E�	^��#G���NT��GP7�L9.1+�C1CF|_�\���W���wߝ[�@TdqM�3S9�������A�F�+H=Uj��STM�E��t%��Ub_��`FE^�j^��ʱ~Wῢ_o�K������HcnE'Xd.�ã63W咳��ߙ�H�j��ɫ����N>�؇� Lɍ�?U��-��ۨp��[��0SL^V:̅w��OG��H����O�)O�,����}Ѻk�x� �
�B���Y�D�um�`�5\Ѵ��ULS��� �v���S��Vp$�oz�0���9�$2|=�,�_���9�r*X�_�S����y��A>�&�K �}@�Z�~�&c���d��yۮGq�PO`�� HU%��'q��a���"�H��b��z� �S:���ؗ�={zF2rZ�R?|���޵?Ҡt#����%��2`'NM؇>�1�[+q�r)ҳ��xj70�HNq���8�����kg2�S�]�W�-�ʧOg�*F�`۳^�zV���ز����L�X���l�b�\�X��Y�~]�y&n��CG\H�2m�~�r�����Gg��I�+���f+V(f����>� �o�^8ǅ��Ӷ�SǬ7PX0��N=��<}�X-x�j^㪻���ȩr{�4�$��M�et]�0�|��G�A������w<'�Y��H���� 8��n�B�N˶|�����/��҃8�T��� hUg�⫵���	��ˮ
U�9E^E���[n����҅#��������Kw,踆��ګ���^��<�)pn?CŇ��87^FJO�2>�q�t#́��S�/�#|�68j�����ÐPQ��������V'�g�M��Zu`>�P�j+8w��}�R/8�\��G%�u�!���2��G<@�j�1[Y<�kE)׃bf���E6��l�+J��7��g��/�������lm�-8�7�!�O��v�~}�T(	��8(���]Ps��AҎR�"�Ry�ί�"�Bvn��e���v�ѱ����63q�]ڊpڠ�����v��1�7Z��o!.��OC�~��2t}*����L�I$����jCҴ]�wޙ	^X��)e�T�3p����%Av��AoX���sX�@5�a�"`��w�ݟ�����?T��^���G��H��X�R��<� U ��Dv��Ӵh-�����xq����+����Z9�^.e��ю�9/�(��p��XYO��� F�������U�G��������>+���Ӿ@�(�;�V���W\��Ä�����{<��޻��yH�����Ԟ��:��'�Q�S�*�p�c��\�dd�^������	њ��K����6�zԖ���۷�'?���O�J�E�+���,���jv&�h�������~�� F��ќsvy�x���#v|�DX(4np��J����-"aQ�pN8��eC�Ñ�/���,n�w~<�!.~�������� G=��D�),�!/(��5��Y���<DV���])"Y�b��wxM���f��*૶�i���֑��hX�Bܣ[�;y�n-�:�Pj�~�]s�e��m�;
�v���ܲek�˷#)�"B1#���6��R��ѭr�s��
��`+3Ii���]��ee�n��Y�������;^���	�j4Ȣ[�n�]{�u��ؾ��/�}��i���a�I���^�{D��۞�^�^Y\���ӮZ�?3;ִ=t؎�<�^��Uk���>P# �����0H��{���ܕ�7X��>��O{���:�&���`��Z��ێa,��R��������U�"�x'+Z���w� �W��I.�b"K-��z�<e�S���^N�x^��d�H����~��7k�կ~�c�<?�J��@a�b�s^�5�)PSz֥:�!�H�T�#�X ����Z���Utυ,.E@�F���9׀' ,�aD��9�3V��?�)�Mk�i�,CZ�Qw�(f����Ms���l�����٘v��z��s��@�o�{,��(OJ��w-S������x�N瀋��	o�>�Т�
^��V�U\�ƾ��_��_��m0����U�7sYr���z����.��U�9v�O�S'�z���������}�P 2<4jW^y��t�-62�<�Ղ=�Y��Ŋ++���@Ѝ�����@�
�Op�~}���h�z�С����o�ӥz�A�"��l�s��^���^@7���\�;��3�"DbKq?��lY{jB�TF��.E����xr��M��`�eRk{��g�D	M��q8���{�oe舁�2(�3����Ӆ;B
c��Y�<w�8�a�C���j_P�b�NF� �C���"@�F
�O<asF��c��I����7�r�l�!Q�_��p��o���N���Vl��Q+6P�ᆗU�
h��Uʶ�.{�*k�>�2��̝���E����a�L��=�;�p�a�^{������g�|����m;l����-ۂ2\m������c�֌�ٛg����Ӈ��z�_����ş?��˯�ʞq�Mv��^���G�O���/�q�gT�6�d'�����^��9��%�@)da��*'X�����������{(ɮ�\x�[�s����F3#�r@�H��g�c��f9��᷍��l�1^^��<�m9'EF9k�&O��t��|���s�ۧk���i�3u��=]U7�{Ύ��6�<����je���Mo���IY�Rs�̝�d͊3L�U��et�������?�	xu1Sis Kt����o���`�ca�} 3ȹBW�
�=?�%�aB_�(���H�Q�.J���C"B�j@��ר0� A�
���8����y��F
! ��~���8g2?���*��_+}q]8<R�EeP0`�1��4X�^�O�Z ��������Bޜ\���n��f�sޠB�O-�N#tC���4��L�RN8�@�2U7b8�f!N8-�\G�n�e���O�s�(;�C�w0�Z{ը&O=��<��C�k�.��^�z@
ټK#r�����]���x�,Y�'���Q�������cn<Щ/��z�����JcґO�����X���e|b�P4�5K�Y�bqT���?��O��x���C��&�Nc��R��8L��$�Fֱk��X��C�����=%�܀���C��<��~�;9�6�ɪ%G�`4�^,�-@lѕ�H�
g
v'�5���k������=7�	�P1���;`�d!a���I��*]��� ���� � X��
�TL��H����9�]<�&X�P$x���964�EL����E�Dx��H 7���Nd,�b�sa����f��`դ�W�y�j�G����Xo{:�^'}�+͍���l\�Z�5V����`�5,6�D5�>�A�HO�ׅ(����6��R�A��1��wE��j�T+#�����HWg�Tj�תқM�T�.G����?�o򋷾NV�� �V�4E�o߷�Y�/£�4������4�X2`M���әH|�ټI'z�2ٻ���.�0g� d�'&�TQDr�h�/49�%,X���〛qO,v4u�{���bs���l� �U�������\WW��s]R�M��A�KJ�c�D8�U�E
n��K�5
8�t� ���%*��%� �c��AE�nPldN`C7��P�q~���a�@���j@b�x6pg��W<8'�)�>1�sM�"�����H$*$|��̑����)�	�m�b�i�G^S��Ϫ�*�CU��Ra�,{x��}Kep`��������S*X��Bz#n����Z+Y̽\.�1\�=z�GO ����U��ɸn|�P�z�>���^�v�^GE&ը�zGw��G��d�X�cE�_��l���39s�F��{���q-�)/�-�6��BQ+�V�IOW�.��F��$��QT+n�Z����,��`��,-kzՄ!����P:q�:��Z�܍ՔH����w�i�6�&Zp�4'�[J�$"��jm*!��u����ez�hm�|,a��.X��Wb����,m5�^ ������sI�8�/x��$�&�V3>%�����B4�����}�vZ�Q�!��i���W,�����J�|�FXc^ ����������a(�C�^=6��v|� �C�^j��](��ߧ7�VZ��Ĥ|�d�����T��	|��޺�e+�������·�#�x1w0���IÍgxp�n��s�:�3���ۗx�&9
������y�]�s���M�����c�V�ϼ��Z�S_��3�< &���C����
�:�L6�`�@b�V�,Zj�<>�)��vx����}���l������©N[s��UX�P�\-
�x�FT�D0
x:���E��~*0�7��ix�e��!Y,~��7(YI�CқL�m�ϳ;��v p��b!+�ɷ��h,�:E��!Zm��S��}�����>R�gx\��a ���&�}( �����8��7�zQ��(�ώv��U%1X��~�a{���G 
��f�}	�j��`�խ�5�=��-�S�խiz�܂��
����rV��� k^@���?�cy�[�j�-6�G.�=(?��֮6��e8�
:�!
J.�1T!
��+�*Γ���Ge��{�
��x)����@��#)W���V���|.)�w�>��^�x`���QmG��.'����Q�X9ࡀ��ݿ�8���˧��8>��J"[�#��ȡ]r����EK��j��Er
��"RQ��"�T�z��p�� ��A����	D�A��ˎ�c���T���2�7x>��b<|�B����]�Uxn�,~"�$�'����r�}?Nx����Yx�n�v�f  �K����
}	��N!\#'z�8P>���:������nB����?C��D�W*��K��uOEe��2���C��t�%|����6�~$�VUϿZ	�=��S��;�}�{���pohbO����"e�'=8���f;���T���CϛM �$��>�1'�*�(F�FOθ�f1���9�S^��4s��ɴn�j��X��8��o&r\aUh��x�u]p��@�,����x��K�\p@䰘QJ�67-Y=����=\5i�8�o�^ߤdԺ��"g��8H�X}GӖ�v�K`���0g1�5v\�\�>�*?XC��;=dȇ������=IZ�P\|nx�a�@��eX��C�/��&(4d�� � ���%+������u�p�����Q�Qt�B�v֔�|w�}��
��q���ճ���o��8��)����Uu	t�E"jm�z_wv�˹[/�J��*�T���O��_�.)���@٤Ru?���½c�c[%naZ~���?�01o].�V��~	5��ať*R*oV�[#Se��Z/����i��~�m�w�AV7+~���~�*[�H���'�L�w�v�Ly)tvYy�Χ��2v��i�+҈��G������w�y���w��][����f� !� �a��tv�?2�o�BKf�4�Ua��EO��?��B\x8����Z����`����2QeT�~�C>�>�n��,ߘr�J�g���b�����Ig@4
�:�g�BKPX�;P�q����hL��a�T�����60M�F�9i�wS��EE �z&e�8�9���U'`1���H�m=2�����,�G  ȥ ��#���!�t�2Y�j��Ke5�ft�ܪ��7�vmM���5�\��A�H��}�z !^.��������X��v���-MUd��{e�sd|�\x����'d|�l�7����V������(H\��7�� ����E ��<������q`M����z�굌��ş�2z��1�4T�hp]�J.Hjűw�q�.o6\u�<|�zX�،p����I\��'6:��yv����ρ
�O��sD��B���0D����������v[�x�X,#�^*��|����W��(8*&�휺�p����w��@���>�)�V(BDØ�g�ٱږl��
���˩�V��=�#vC�����C���0%z(#B��q���l+a��6{`I�Ž!���G>��%�5p�}�c�R��m�](���P�ꀾ� �Ī�e�Y��[&�;�-�$j	�=���
��?�8����s���A6�K�bz?�C���iY�f����*��2tx���&&F�d,�.Hhn�z��u��$<?b�L�b��� ��͞������&]w, +��?�����~N]��y�.�$��8Ir��K�\i�yZCjX�ӷ1/�5�����p�c�(6g5j;����$.��a�ǯ�3���%a>O˟�B�,c�8�6"餱|��iE`�g
��(?���{���!A���Y?�����-�F/�`���U}�X=�%r�Tn�}p�O�Tq����L�#\w�QC�� �_��_J��0ҡ�$l֧� 4��u���Kj��a��AȝBΘ�׆36�5��h�ò����C�䓻��-���Fr�q���uq��>�e3/�FY��? _����u��U�rM]���iG<p׮r��ak�GͰ^��Ns)�q�C��p<��|�3�7�Ɋd �#�V�+^�
��W�l^+�i]�ӗO�v|R'��dCv=�CjU��֝��@>+�5���E-�T:�����Xp+�%��'(F�W�p�P���'��yQ��µ6����0"�Ճ9gXe����e2lCd�X��7C/[�Z�:��q|&*B;1��҇g�d-�E ���Bx#�okk�81i��By��l��R@�*Ž�F�#m\�į �݃Ec#�q���ڄd<�1�E:e׳~
4϶XQ��������A��0�BD(��Ї>��ϸ�gp�DZ]�{�!�6�����J]��d��@�����<8j�����l�v�z,��� %�m�}�d��5�i(x�q��V#p�bb�(����N)td�%/y��k9Ier�eW�Y��&IN6��*�U�����1w�?�c8tP����ֹ���k���H�R�����k������X��Q���]ۤ�_j�Ѓw�#�X*�:�gƅ��J@%�d�.�?�.�@�a�<����r���ܡ��pNl �5躓��վ�L����7��S����?���~׬Z]S�@y& Q�=6z̅�j�%䦳7ʅl3c�;`�j(�񊅐�� &�>rԎ�Y�0�rd�����{l=�
7(�8��EBki��a����V����P 𤡸 ��}�8�����Xƫ�Є�f��ի��[��FR>�����è��F�[^�R�3%5�r�K�������ռ�`<��/���y9�c�~�<����84��+��I.[-����\�(�~��!�c`rtJ>����C�<x\�x�(l���s�J���}�0�x0�L���p��T&�~��񉒹��t`�@�����pb�@� ɋ��x<,�~c��*!��.#,�|v&_���6���ŴI7hd! @��
S
�C���,,*�zc���D�c���  �ň\Y+`�!,�{D����m�/n�ه�an���<��>{H�;M�	�i�3��:,rҋ�w�e��_�m�ug�  q���7|���Hр�`]�<�'�>�{"�k�9(!��\ӣ���v`|8+W,�m�oAה��!�`�aF&U�wu�[���j7xwu0���$���ɸ�g쇛~��O~��	����J���M@�Q �	��,�[�J���$U,tv�cO<n��@A��!_0׋Aӝ��?��e؇}E��"��K�я~Ԅ?�
؜�dY��H� Ə���b3zǬ>,�?��?�ςW�f�|�4��bq�����gB��⛵:�B�T�'Tk	-��h�`Ψ�Q��m��CH���j���.�s/ ,0Z��� H�`�ạ�|b7Ɗ�����i|ZgZ�0&��� 7���7�O饢0	��[�����ǏkA��A��w�wm���_��	i6H��>��4��:X5�A�c���뿶�!��ϡ�PQ;T���&[�c���9���i�5b�sd^���p*�^�Z������\���s��z�"�^�|Y�|�]���S���j�Q����|����8��q����D����d��/����b��)/��d#$d.2�Ҙ`,>L>�U0�c��7,J��ȊȒo�ƳM#�}>�O��C�~��`�����;?��D]E��=$��b�r�@#�nD�"����C��Q5��mm9���h%B�����_h����{��d
d��j���XD^��/��`g)���>�|����h���a�\ ��{�]���a,����`������8'�C�<�������ll�C>�=7�R�,�FՅ�@��ϲ�{�T�޾���⹌�=��F	��� �R�*ܔz���?���9E�0����������=<G(W��^ �'�7�1�02�9������:��|�5~r��˰i�4�7��eec���Y���������0��I��k0�E�&�	�釞����EuH�<��s��0���Ca�L���U��2��m�ԋ��&|��ZG�o������m����Hos�~��o�+��aeb�A�����p,��/�.,�w��]	���!�������c���#$�Bˇz�ӦWɦG����i���<����M���Y=�U�@���7��ֿg���۴Y���K��[R���*�S���64�JK-UK���~��Y�HH�sG�������C���O����-���bIVi3�@�EzrW ��S^��7�Z�/Fg��������d�9��O���,6,�>�$P��d �Gr�%����o��L��:J�;��뒎�ZS�qݼ�p�k�}#���:�7��!��	��[�J ���Φ����>.��8�AC�\�X#C2n����7���a"EaϺV���%��3Ɍc5�c��B�'`�1@t�F�*����A�ǳR����'���w�Q��f?3�Dm�r��V�4�����m�:�+ӎ�>�0}d���������w[��Ph��½HXã�L���C��DC
���3f(��c���c��b�i/�1�L\{̰�9>���
�Ho��\�x�X�
��P ���U���[� V5?ϟ�l��l}���oTC)N�%�B��KnNʕI��fBG�4R�ؑ�ſӨ��F����n��D-�b!j��LaDWߧh�����rV���X}�(r�P �*��q\*,����J���P��	M�@������@1�G\��J��%��ҟ�]7Ce� <�??�R肇�ew��fA��y�汦,\j�9�_��P��q��=�1�"(?�opݸ�}�c���7�5��"�3�O���lY$��>�~=A+l�?N_��<��R�\Z�\d~۷Z���9c�<-��H�!��W.x,j|�)3�˦|�87,�Z�YS�	� ��e�?��q�wa'�L�l���j(�0� �AT!�,F�i9?l��>e,�n?&;�:k��(��!�?��}( h�0�DCk�	��6\��!b�T4P��nR�!1��3�l��ռG�Q��8��CD>�r����Hv�V���!��c�L�d��P8a���֫�7���q�?�9~��=����?��$J���L`ؓρ�<�$������<��fΆ������Nߘ�|�_�>'6�o��	�kCDxDJPX�'j  �a ���[@̵i�$�oq̮�&�՛����~�)�nE
9wO�c��6E��[D���,��FvōG+�����s��%�[t�3n���R{,l�����/���6��/0(�0����g���}�LBC�x��|H?��?�Z�~�����ѐ	F�/s]��ܵ.\�а��Z��n�\V�"0@�{F�����2�t�q�)��2K��h�^)ǐ�ؓͪ�E�\<Yw]4����	��g��)�i(����7&������':N{����;���VN�oՐۃ
�V�����	��l��e�p� I?"�=�S��Q� ��PO���ftb�^�D�T���F����9c���;�q2G�e��o�QPxFC̅w�1��\���;(MT�T��F���#�?$�HoϠ�^�A�U5�O(N��%��f��	z�T�����"bh�ъ��|N�"�@Z�E���IfB&9�,�ހ��i��!Z/P���s����T*�w�voeA7����r��n]��DTܗ���V��Cf�l����� �Q7��@7�Q6��+Z~�M{<W��kQ-q���ټL�F����K��ua�Fv���9cI^�74tHB$��h�3�O�"�3iT��4ʡ�-�8��a蘈?�C3ĕ��Ӝ�8��|��ӧn�`�#Q+��LK����f��|r�3yǇ��{<�}����ύ�$�,����T&[z�r�H9��(t��
c��b@Ӏ|�]}�cm��8�cv#��]����n���o88rW�Z:���V�e]]0ҜYŔ�4 %p�l���}�*x��"F߈�	^�b�:��̣�8i���"=�٨���4����  ޘ-.��Td8�w�h��°-v��|<.CA�|~a?��\�KK�_�R�ԪGb\+Y �b��Ѐ�Ti��LUʒ�,>ZE�_��u� �'���Ӷ���6f�I��v�t���)[S&4a�u>U�X�s���|Q[H��ܴ�vh��˷�����'8� �a�Ic�0�I �oȠtj�{��TP �L�_?Q�[��<O'2Ny�?''r<U���3���	.�����Xt�(�}aތv���Wr0���#�J�xD��k�f\%��
�TC,�+99U�kba������7Bc\�f��Ԙl&������h��5Z�HrhX�rprj�5H䆇G��Iވ���d�*Z.�^�W\_$v��'KR����d&�l͠��p�&�g�f�0����~Q��_X���F���?�8��f��%N�D
pChd�3�A�؊�������a�M<N
O�]��Dt��&u����bh)���D[��{��T,�F(�uߨ98_�~�]����I4��26Q�#G'��k��ϿVV�X�\/��M��'{�Ʊ1�T��w:�����ό�J��zcK]��K�O�I�Z3�P+�Z�
��:T�ҥY�'P�����U2Ĝ+:K��x���]�`}�^����V�Npq�fU��F�m˿����� T��1�6�\�p��er��73X��&�7M����y��կqpb��)Q�ҝcl��u�`Xv�6�Å!:ؔ��y����ʰD�8��1��;��T2k��U��C����%/�ŘH��5��7�~'�W�q<܁Mb���dE��>�d!�	��A�h��Ȯ��Lޗ��I1P�g�t�������6湟�;��u����毙�ol�56wMM�y�Ӵ���<���6&*����<�Y�ef/^����Le�4,z��Ҥ|���_��~/e��W�6?�/��[�o�Z1A福u?�@��1�f(�����8P��`�.�#�����d�gZ!�o�:����ϒ+.�\���oX%1��(�:����x�Є�iZ] ������U����'�z����1{9�r �=}�d`�Y��=�׼V�{�L	�(+��u�Ԫ�U���#�
�Ը�FG��L�wMi�Fdx��f#2%e���;W�V��b���d�X��K�����G��^3���
�f:���2��%�Gk@@4*��<���(x;���T��3�!�V�7{���ǧ�f3�ڨV�,�0��,��V�..�!"q>���n�.m>%g^Ohg�3FH�7�����$��$�%J�e�&��I��H�V^q򨤲*X¼Y��;0��E�S.H�����y�����y�E�P�J�)r�/Z���@��@?�D=Bz@�`/�3�Z�l\n&�c�PF?�FG9mI}�&�׆�J@�����u��<Fz��?�����"_E�������Ƌ��c J�JY3p��L��z,E��V�?,GF�4b��.3�4�'��(X����Z���L[��D������7��g2Xc�$��|�͇tC	ԬaRl��=i^X3���X�˰k!�]������(��aPV6tx�>�d�R��R��Ȧ�Ζ�k�[�� ��ߡ1�N�E��E^QԂ��r�
\;����*��ꄏZ��O���k�����I���/�X�ٲU��XeM���j�`e� �h�fO,�׽�u��YD���ˇM��D��d�"����0b�ȬE�o�,��}��45i:������czh>��kL�h�!�'%&TL(�@d�d:�_u�?2��@������4Bm���7��u��b�/�G7r���w�h/��y����HP��JkB�}&��#'\U���&�èG@��g2ܚm4 �.���\�}P3u`-��}���~?��*��ç�-���	BrhP
�j�|̏��X�7l��Q�h��dVn΄P�2���Ϫ������ร�_��-�E�Е+_M�=�x��GT���8~E�F�u0.�鄷	^���GS�h�X�O+Q*��8�c��T��p����}g�/���(�}�1t�1�U����T'z0'&N����ȇE�?�}��(䬝㱣#*�'�|\�������q�9r�ŗ��3j����?޾=!������u:7po阡�I� [��u�\�|��pJr�H���%w��=����K�汪�h�����^����L}@Xl7�|�qsӊ�5 �>r�B�;���<����_�z����[,c�� oj�+����Mق���"I�b¬h4��E����&������|�=��A��t#����ZY��U�(̙�`a3��1��V]qI�zL��n8P��YG��7h՗a�=4�?	��x�e���sq3�,��~���5,����F�	�Oڊ�,~��±��	Ⱖ�جi"OƦ/tmQ���҈��A6gE;
�nK����������R��G�� U�j���5m�tʅ$Cԩ��~=����P�t��$���g�W�<AJ�����v���,O^#�a���$�3��E�Y�<f��;N83��0%Qz����Y�C���k�5FS�����@oP���������߃�����7!{�<!�|ر�I+P��p�9,O��>����] ��Ke͚U�8��'w<������I�)/�[�}�[M��<O7�9��f�c�%���[�˭��"F8:<l�����_Z���{�g�a���2��6l��.���P�o����Qs�����o���a���d%8O���>� ��:�ıZ`Q�*�'�N�B�gI�,�����QF�$�Z��W��I��.����P�V���<��*��n�JY��B��9"ׂ̡�G+�!�{� �Z��j2�|H�S�:�[��j}DJ�q��(�5e���;oT��Vc�!��]X�8_Ը�(;u�"�%�!�jჷV�U��KO�R����E�*m��N��`mG�0�9*�ָ�U^�q�:�*@Gꗊ��Gus#�l�r΀���V%�����U3�d�ff
�|>Ãa��-�Vፐ_:t�j�ٺ9NVV��6���
��e�u��ީVc~��ǯWFr-�����Y��>��"��L�����`���"��_��������@��=����j܌���!��I]�����3��(�՛�*���-�7��笁;d���0W��
~�S^�����q�s&��͛�ڄ���ʷ��e�ֳ�uk����	�6fdl|B����	�y�u�]g� x�Gy$�h�F̎�V�h,�p��2f�����2�(�}S*�U�,D"�j�J�B4�=I�f�E+{���M��5 �j:���F�4�.<�r���g�/��Jy��+׮P!1�B<vC�p^�:@���ty�*���q����խ���C~�
��� E{��321Z6�epi���,Q-���+��v=.���p�K�8�B;+K���a�H��UUL��0p���T,)it˝j�g����#�^�#�s�'���/�;������REcޢ�wthJ���άtvAY�1<�I��g6�#E}��[��u�ͥ��)�� ϰ&��f&k��,��nTu9z����O�9<t����N��~,������cR���r>��I{,�1`U}cF�k_l����8b.�Ǽ�����n�[ �B���z�{�k�;�������=�\�T����񈮑��Y�D��)kh?Uv��K��������;�'+V���/���m�'���>�ih�e�<兿��� ���U�;�Q�������q:\(&�l-�p��B�S-�1k�v�-��%�Nm�����	�^ U��݋�/��/��@7%߭$wG3�ۉ�f:�f��E��I�m�ΕMg�։�������*�.�_7�V��@U��C�F�;������b�'��R#�.�ۈ�#uRy+V{��G��w���뮽J��ҮQ7�5��Z�D�#�������wn����u�Y�e�:U&�di����*��>V�o�^��(ʍ�]%}��t�۰�W#���kBqa�'Z&Ǝɒ%r��W�v^ ���\�>�HY�ꍤ��Bjt����#�ߴ������*.T���W���[=� �8�s5>V�o|�G��^p��?�i�/��!��IC�c�׳����m�,W^u���Y�9���	�F��R1���}Xʓr��[d��:?u����[�}ʱ��7��GF�^���K����<��E�����0���V��O2|�B�������~�+v.th����Д �������#r9C�航���xTe�r�?��q:R��2/}�K���蓣:Gw��r�%W�~h�ʕ�������f$���k1Ny�ߒ�'r�-Xh��Uj�8p�ڿ�P��֩��::T"n��*�qO
ZZ"����H%
��;�y�?��/ؿ	�d���\�6�
�|/c�O3���#maX)(�)�&�,*��zք�6>Si | lr����VQ��ch��k��"��Q�o���@Za������MB�%��e�S1���ʢ�	ز*�@/���`��-��p�f�︡�
�M)XE����q��B!{p���Y�5w��]C e@��oOA����Gz�s"��a�,C�j��u�A��~�
���B��Tծ6�BөF$��6�8!�Qu�"2�IxO�������Kh�fG��(���e3h2��zQY��	bNcsGx����p�0����@	�z���Hf��q��b�q3RH���kD������F$�eMJ6������L( �u���
�9��!t!C�^�7 �@����/����jҮbxl|D��R}�i[��a��	�$��󙔮�kk�DgGo���:�q����o;�����Y��h��8D���ߑ�!>��x8��@1��o�����P2l���|/����Ic4[K��ɒd�ŵk�yF9�؂��'"5WSV6m(���+"6mEh%�w ��<F�v�C@�@�{�X]��Z��[,��>+��Q$�1��	,$N+�)��ͨ�"1�#�آ�N@:�G�a��į��\�ؘ�rQ�6*��UХ$��}�*$�E*v�Z�b�]U,���M�EU�����nT$V 4K����ҁU7!�S��͍����`���K��T�~�
�|���ME�Y�Q�nM|`������*�lƞc��C��)�C�-}h�':ȕJS�iK�?_���3H�\�F�"�i�0��.Yh{*c���ײ�D�I�;K�B'��b�'
}�A`�{�{����ޒ��?��^�*���lﳾ�͎X=��Z2��^!��kA-i�$���&��,��`^\�:��n�2��3P�Tͪ&�R)���>�.�	F��	���v+�5	:eCnQb��+-g%=<�^z������7-.�������/}�K���`˾���}�9Z:���9�9Z)��,�kp/q�˨��E��*��:W�Ѕ�`� �Ě���3b��#��Аad �g"V["^\6��x,���5�Q�)�@b��0F��s�H��0��$���g�TW��6��nө72U���В�����d�D���x��A�ϪL��.�	(�sʚ�l?D筼���E�(��'	q�!Y=^�����2錛�c*劕j��	{�~Y�5m	_�S�u��z�����\C)�)���=8�qEP�_#w�$�[�<s-�~�O��a�Cj��:m�P�r�����Fw�>!�Hp߰�Br�gfM��c�Ν������oΫ����q���8�RdH�l��F�*U5�
�NWcr``�<f����=.'�E?����?�@U`GgA�����Kz�j���V�[�{���Y#���L��DE��V����6����^ ,�������K��+���|�#����\@$��U�ܠz�6}͌��۳5��������B�)uOIU���`�Y*X�CG�&�!���F"��F�j9v���\�g �[�`�a�NQ֡�fE̽��N����D�����>��g��ʆH*������g����1�u�������]����%a������5�Vv���W��UG��r�p��BcYU�cG�z�D/�`�����16Z���^��;t�����|%e-���hk�3��8����
Wmj�Gz�X��$�#g)�JU+�����̑#Cv{� B38�SQ������U��l~�z-׀�9S^z�\u�T&&;,��/��B������wK?��Sjh��W�hG�L�2#'��ǖ�+����q��gn=�Ċ�0�^��D w��;��p��� ��?k�~���uk7ȡ�g���V�����n���~����I)�|��[^���zpL'ͫX�8�$�%aN��54я�s�v��7�+�-W_�y��{���.��]�K,|�u�u�M[Wv�aX�F�W낯�ӟ����P7�t���o���0�~s�"7�$�o��o���E鉺-� p���b���˖���:Y�|�)��v>)�?-S��%E��EY+r��`�2Y�~��%�?�^FT��ԣ���c,�L�
�^������;e��5�v��1cC>�o�ZS%#��d:,�X�5 �*��'�fQ-[�Tϻ֊���{Z���%�)�\R9C� {_l7��8,��@��߰BV�Z/�� ���'ǆ����,T�kjD����������2A�D歹�T �-Y�v>*��~R�"ٲ%�%U�L>�)� B�%�ӻB֯9[ϻN��1����U>�T����K>�ڂ�)���\��Ⱥ���Ы����?�C�ј���p���R4�����}:��e�ʵ����d����Ԩ	�P�	sVL('t��Pa?�B�]+T���9����^��\6{MHDW��؈��4k�DӍ��j�}�8��1�.��ϱc�~��_��_���E�@����Rٹ�aٷ��Շt��V+��;��e��~y��'u�����,�F��@~ͼQim�EQx��}��#
m��bR�㮻�˥_&�j�#q�~�9rdhL���'�ʭ�1n�p�W˦�ےb�{��\>Ұ����`�����|�k_��Sf��1��s5��q�-�GN|D�C=!6�I�Z�Thde�곥�g�
�N�9��aCڬ��#G��sm�����L�����9c�f�����W�궚
c��Cf����X��D��2��@ϹV֮ۨ�YH�3Ղ�{߯
V��%��q�����w��sW��X-����JU��U9��rŹ�, ��^��N���M�.TA![P�Vz�d�؈^g�u���oZYU+W�wْ�r��3�"�ϓ�*��� @�*F��Qv�O*g�w����z7���*A���;/��R�Z������Wb�@1V��~�w�Z�)Y��G�?'?�~�
"�ʺ�v�zC׬�?��/���v�U��4 1ͫE�~c�����x<nq��-8�A� }Fh�۷\�:{�z =�,;{d�*���wD�1m��P�5Pn4�T��I����ǯ�hQ+Xf���]�z�z���~�����Χ���5�y�����}�3 ��[���!� $���սT���(���W	dr��Tv��~�U��s�7�h�Ȱ
�$\dJ��1:s�Q�Mҭ��#�������E/ԍ���^)W\q�Z~=�l���[�����.6K�/~�f���H�7��|�r�ԧ>eP:|�w~�w���a[��,�&�n!h.6���.���A�U�ꆯ��4fbq�n������.��YQV�ZŹ��~��4\��b��,��IIO�r�n�ֈɺ ��(O��c!�jC�Z�pܜ�TEܻ_��B-�^�2��M�b�UƻU��ˤ����T������Wk+��2���:u�;:���c&�sªY��l�*1�x����kM�@L��V]�� ����4mJ�����0�TC�W��֯�"#c���ڛD�4��F̀M���):O%��"�*�^�R\����H�`���z�=�dD�j�58�ӈg;Σ�s��J��Y��jYv�K�=�d�>��S%QO�1�U�T�w}E.o��z���Md�h�=�R�3�@�!��3:��~���X�L�
�Azy��y��F��Ac���%�F��<�P"�x��<�b�WR��q��Ss�2,tp}϶��ׂ�IՀC�����?���z��PBr�礝��<~Ȋ׼���[��,]��y���}�?�Ò����r�5�ɖsϓ��X���>�_�)����e�����?j%�<��U�� G�O"����)/��Fc�V���kn0aE�Sk'�ﰅ`t�z� �	d�X�@�� �9T��;��~�#y���-+W��!@iU,􁲦�O�2>Y_��X��<��,�zF^���e_'�ͤU�Bh�^��
��7�u����׾c������j��q�*���U2e�6�I�KRQ����m��yz�nٳg�\r�r����E��`�U`���{���&J�Id�����˱�1y�^��?_�EQ�mJ��
�@�W��MDQά�~���^��]�����ea�[o�U�٣Ϸd��(*������yq��n9g�6����S;���[/���&Y�r�Z��l��.[c��)��`�U��7�\6o�P��|�;ߖ��k����s6� �2B2��&�`EYl��h�֨�c�paC��?���ۥ�җ�D��id�t�B����*r5j��]{�z]c��#����9�\ 7��")輢�"�Ϲϫ�����R]��.ٲ�K�~�K_�b��oy�іXD�i��_��z��]��D�r	�^Bk�C?�ӞY��î}&@�R ,�\�
}�pѡ�:��S����ȵE��>X`����@fpO���� Q���A��k��P���s�̳Αo�9�������iN��d�$w�u��w�vɫq�~�1��g�o��=MNy�H+Ӡ�����y)����|�2Zg�;� �����N��z��g�����.��� ��g�/$w�	�C�ŀ�x�Ï>��lC�a,Z�-��8��%��	�@����Y#֟c��� �DW�j9��F������r>2<)˗ʹ[/�u�W� ,��ZX�g���Q��t�jA����19phH��v�
��,TS�ؽ
�2b��4�,H��D5�9����e�X��.�B�ظV��}��rV��87��0��eЩ2��Uo�wTWJ�l��X��b �ƘP:��0|Y��2}�y��'Գ�+�ܢ�|�����Vv=�A�!��"Jg����S�6WeAP6��@t��X�X(-g�EC(�]w�t� -�>�J����BY��K�QŠ�H2#4�0�Td��U�۷B��T{r���?d��\v��5�B���<G�0���e��Y�"/G����[^�U6��Y�*�.�Y�8�"��!��ݳD�Z�z+Crtx��vδyH�a�#w���q�.V�������9�p�ؓd�D�Ίeˍ��!_|�W0 �
�0��rYX���W\j�H��;�����s��##���ʑo盦T��;t�M�1WP˜^��K�<�pp������Mem~��ߕG}��;V�Yia��jo�;'���wВ�۷ߗ^r{�!0v��8>��Z%0*{�0�)|�S�4�Pr瓆�ս�	o��<���j���f�	*#n�r	N��']B�^u�!�9���㐁�$2N]-�RmqC�����@,�6�Ej�Ud�h+��JĪw+�X!mU�)K�A0cn�F;²�LNLY���c��ڋ�W����jgü�[��l�f��A�r��>���9���}��҃Ŗ
�"oČ��Ɋ	U��1cNZ�8�\6o���*5�r&x�:�]�H#�� �',i��@11��h��C�P!]��˲���c�5㺪��X>��Ƚ�T� }�g4:6ay�FX����n(��Q���x��F07C��y��F�,�B��R��ks�deGGg�9|�L~(R��=:iV�Ɛ�(YL������>"�"�P��8�~�Ϳjt ���� �9�����Y�c�+�
|�+_��M�e��.Dɶ�!Tv�ܽ��ͷ�q��ۿ�h��ET*1P�1�ZgA�����.�
���"&��V t��
�q��׿f�<�:� �U����x����ZR�0��i�� Uox������k֭�߻ݒ>��� �/��/m��B�G�����E<F��b�%����͊�@�WtE7i��8��u��L�"���$q²��nk�ё�!�mxR;G�GIP���0�՚��;��B](	�x�{n}"ǜ�U�?.	Cᙕ�QRp���¸f�Op^��
N��������g�{�.�7N�ȑU�K7�y+�r��(�M�TP�������I�0ra���Ūa]���)?\c*��Z��t�
�i�hV��P˭jJ7g�s�X�*�1Q��-����F��rE]��F��%��I$K5tךN�cZr��A �2����m�y_4��i����Z��>L�r?��e@=�?~ߟ�
X7d�>�Ʒ�������>A`㻀h�3�l��`�=�z]�o4��5BX00-�{�-	�#g\�l�m�>�[��X��c�R?RO,k��uu��B��[�(�B��׿�����`0"��'4>ڴ�9��2��2�4����a���&�1�npΨ� 4��̊h#$R��>.�g2nz��������n.X_��������/����!��^ ��@k�����2I�)�K$�`(���>��D">����2τ���["�P�g�OX��ݜ�*DQҎtnn)Zˁ	m�1 �,����"b6�~^㣅���ʙ�U�m��3�<S>������ߟ�� ���>�9�� ���D�^Ƴd�ܽ#�����T8'�|8h���s��6��aʹˎ!�3��Ȋ���ݴX	�B> E]�Ї�w����躄M'pY��\W���~�17]�t�O{ܪ�Y84�No|&:_���{Z��k��5$>����54�H�s��b�3���b�}2�{籉�'j�J���G�h���量>�-��AZp&�G�b�mmb�B�`O=�>��>�k����}�'��Z�v�F�욟04��W's�s�<�,��:�+rv�x ��>�,9�0|zOT4Xg8����|��8�k>�|�M��40��P���zh�aa�+`����O��L�=Sc�{&i-S�(Y��s�P8aP���rS(���>-5�"�{���M���~��;�w)l}�#T���y|AO��S���Ӓ'j������ p��2!Tدi~�|^�5�3�p[H�p<�ab��B��ÿ���.�G>������yoD�  b���-/ �
^��,����Ƃ� ��c����hNFs,�����ɤ7�'�m�i�yc�Vڇ?�a����}�����͍�>������7�s���P��L!�6�/�}�I���'��Mkʷ�\«��"6Z��5҂Ǳ���hnxc��y_�ӛ�s$�Wz$ �W����d(�a)���򇉀�����2���sH͖�o����}�~Z$H�4?,⯋VU긎�DyF~�g���-'k�f��u�w��N^��#��yDU?��y��ו�W�>���4p���q����O�
�h�%��Z9=c��
[�M<<�������>p�xA�#�e�^ ��6|Z�'{���!����+Z0��Z}��D�-�wz�x�gU�|�<���r��js�z|���|___b�3�G�L�B��p���A9Vw����������\�����4�3ŵ���yzE�Z����q�B�
�G����g���O:8�4p0'�(j��Q���ż�Y��+Þ�������9�=��Z�4<V��6�ۉ@�hٙ���Xsq/��/f��_d�6`% �	�I<
��M�\�}ف*e
!*1ߺa��0U4� �.9|d(&�j�X�͞�h���	�5�����c�3���5�y����=2|Ԅ�/����A�{�@b_���{�6L76�o��:g���Ő_�`}߁�"�s�u�b뉰�ߙ��@@�Ч���5%Z����>�(]�������-,��c226*ݽ=��:p�����87���8�x�~���:������>�~�]Ιڢ�c��:��,����Q"�S��[��g�dz���a��k��c��h�y��j��Kn$n�<^�uIRaa�c0AI4r���'�]��� �}�In��7�Ip�����l$b����L�����hY�@K���b��ap�O~�3�r4�f�Oa���.U�B��U���3ă�
!��.`�Y�CagB ���x0����܎�s��)�}t�����ߏ�7���00�Al߾݊S�5@1c#oT��n�5����2����s�d3��*w>_*zz����yP���<=��Ѝ�Ȍ��}���h�Od������ډ��L�Ml��+�u˗��Ń��H��p6)�
y�)q^�8�no��	&?]|�~8p�\�/?�����8�މz&�p�΃��_&�y���jm��9?��G��������ix��G�c���Ƿ���l(��0�
��6p�L��a���OC�
��Nǟ+*Z�;<��;���i�%Iq�A�`��V�)�4�4jq_+6#Qb�"�/�3hm>�� h�Rc��e�_�ͮ��<%]=�I�̚�x�]Za�d`�b�۱�ߌ~���Lt"j��h��76b�� 
����Ď,��~T*�d���;�8���<zܒMq��k1��s�a�#���?b��0����%T�I &�zg耉A?�K���R�;3|�����{)��x�����G��|�|��W�6س� �ņ�Oy�?Ο�/^̔_p�lݺU�����gYSr��!������S;-�%��'>���F�{��x��]���+
�V{��s{�'�g��3�G�{m !g�
D��oȽ�w�}VD�y�o���>Aˬ�ʳٔL��I�?/<���u����љ�Ze������p�g�s�>tD���;��"y���70�1�D�0��dCD����G{�������ʬ{1���g�^�k�J��_h�a�Zy���#i�a`":1��׹�|����i���J!!iֿ8��/|�M8NWwG�Ks! s����@ׯ_/o}�[�c��ii�~���Cdh��t�~���¥����h��h=f#h$z��믗[n���	�@0�g��-[�X��Aw�u�) �*,��Ny�ߘ��
`jr�������w�g�nk��{�N�x�K�ʦ�g�E�\f��(�B�6@�|�I+��
������_~����G�h_}�7�Bb�l��h��6RG4ú적~�K^�dFz{�L^ �������ADa��A��W��UV=��������F���
9�A����W_)��21>"#��r�]w�~U H����DL�<!�<|�zc�o��Tڈ�n��K����J�/}�|�ߴn^����jU�h�N���NȘ��o��h���O�3��W�C���GOW����ܿG����㏘G��R(�#����\x��&Pdx���lE��n�8b���Qs����s�\t�����)�V�etx�H�\����4���l-�j�>����ɫo�o���E\(w�q�'&�T���_ϻ�
��G��*��l;�<y�������޹K����h
 Z��H kBҎ��Vc���^'g�`�͓B}�g��^�23�ц!�B7t���o�Ċ��Rq�%�ʚU��V-�qZ�����cCOKg�*ݝ���RW����DE���w��񆛭��ٛ6�k�<��&�|���*�����o5l�!̢�}��_�ݲ՚z䳁<p�vY��G�ذR���ɤ�Z�i�6���P�~\?[S�������ꪫl1��G��6$�B^�}�{���7�2'�3���e�k��h�>�0靣;���Y�- r0������mo3��=��h�CV`�W+E��أ*+�j .�]�G%�	\߈L��O��ب�i����++V�1�Б����,>�:=Q�S^���a1�C���ի�J�^5�s�S�f������J��Svr������ݵk��t�M�;�Z��v[R��&ޯx�+l� ��\>(P=ca���( j��o��x��3�>��C�7�7I#R����W~�W����}��=],����<��òn�2�~���J:$�=-wv����49w�6k�y�g��e+�����/����-�g�
_8K��T0�)�I�VD[ɻ�O�oe�֤�!�0m�ᒱ*Z�����xa1@�Ӫ���+��������ϟ�V�!IZ{�G{���
\둃��;o������9~�������x����qR�<�{X����+�FJDVƋS�C�\iX��{�Tt�=?�W���Vk�T�K�Z��c!!�S^�A넯�42�M���{�|�;�J�h۵�C[?�'����/ ����/[|n����>=�y�<�$vj'|O�A�.l�9��G���>��gL��;�A�S�oذ��;�������-~~X�4�l�֟�0D���dJ��L8ցj��EǏ���	�5�Ԩ���,j�'lT+K��2����ٙ��֟4���0N�0H'�Ux��ĉ=8Y�����q�Xxn"�?2��]w��C�����0��h��;��Qx���ַ�%��ޝ���T�-oy�y�0����]�ش�'��P�̎�!'��Xod�4ʖOѤ�#�$�I�����r#�N�"�(j͞��4Y���ʥK,�a��R�Eƪ�J�%�q�1�ή��d�>�B�%~H�X����������\>򑏘�G�7�����Ѭ�����sj��>�0�[����~������G�O������˭��j{�`ޛ6m�O}�S�؊�M�H���/�5�֫LI����AQ��v�9I�p�(t��XY�_�m۶%b<f�"?�0[×V�/�a���
�y"�Zk׬R/��}�<�G��0�U��/.�JoO��-H�|P?7 �]v��e�>7
���`����"����=��K��?�qz��m��>(H��=컀����{v�o���MX�$y�������ꔳ��,�G��ɤ�,��υf�����6m��v�BG���	
F�X�q��iKu��R���]x�
�,[�R�ղ<��ӪaG�qG��!眳M.�����I\.6r��~`߁���|�8����wZ���ɇ��}�p�c�N�ʎ��q���W�'���ty��"��$V~GRg�d�YB�0�o�1[���,77)����8?�/�ɉ�K�������y�1�_�2�JƻX�J��5*  ��P�����Hދ����-$}��o �?&79�lbC�z2T2��gHzs�}!�
��_��s0��k�:�iP�����y�@��-��y�_����~��,��<4�1j�������?o�j�$+d�X��{:dO'��U���Y��(%K���_n�Q�����]O���s�}��������XИp<������=G^�����1Y�t�\z�UF�p���Y��T���˖�%����bIg���m�<t1$k':>������ :,AI����ÇfsQ�Q��h�gjpsb�#?q�����E�M�E��^@;�/k�B+�\�>ԕ��A�4�����m�=(x�~c�R}�/R��^�7=�`ǿ��կ���ߟ��=_1P]s�5r�7&�W���3���]���j�H��e/7K���&,2�DA��%�B�G�߉ޢ^7�F"�}#ȓ�o�9i��+<���$i$�U�A�1^�\_��WY���0#�a��?���������{����<�B��������0���<�ɟ���gC �y���׿���{��{6Ǆ{�a"$���"S�c�y��j�wȗ�����K�AC�=��/|�K���_�x��s�]�?\,��2��Φ��*��k}�s��z�^t�ҥ���yW��e�^���JZ5m���9�Q���6&������-��A�nX��n m�o��o�{����I�+���bwl�Mr7�W����!�[C52�%����䴾[?e�9���6L�h8f�7+}�
A:��Z���(�sB/D?\}�����/]�tV�����ph�ؘ���&�9ر> ��}�I���JdO?l7�kn��|A�>�LY�r��3O�^j��W�=��q?I]26���
E%9�u���S��ӛx"~��38z�b�	;�[�͈���k��<P��MG���,������gϊ�J?,��`�����C�����dQ���k��mF���d��+L�A��=��a�!��q�Fy׻ޕFrmq� �eq����TM���׾��\W�<e�RД��)�G~L����q�d��F�q�� ZP�<ɚ���7�pú��߿�v��B]f͆�=�Ѓ��s�w���L���zF�����#�=jud�%���~�*&
'Z|X���o!�b���UNE ���R�c����p�v�s-~��
����ϰJ���ߧ�dώ!!�W�ӨI�~��' �q8�^�{���`������8Y�ʕ��?/�m������}�[��l����=��a/���'�}eϵOO�k�ϖ덞�=Syvqs���uB@c�RI`��'�y*1�}0�_��,��y�fS~��{;�{ts�X)[A����g��/�����i�珌o������RR���f\!&Ъ��/+V�2W�O,���a�����zUd������M��0�?�iq�9n�W������l's����xa��%c�rȑ��^�|���� ^�������}sh�֧��I5X�xQ�Q��q�p��S�u����a�ؼ����xp����1i_����5���=�䥳Ё��f��rQXO�+9j9�T*�sCh3:o���뇑�^D�P�B���g�Y*.��(� �<BZ���%�^�'~�i�|�s��yŋ���/s�}��)=ey���>ԓ��~����7��]?>��}$b��Pq5+J�#��a�֭r�X请�[�T�ܷ�LV��l��~y����D��Z�I6?�C�NS���rv�:��\�!~%� ���?����d`�	',V$��.C01���OǌX���f��}�!x�,xp����7[�>� ��O@���͍͌P�� �i����`��%�������7==)��5��7�,T
LB#���~7���$)^V^��ot|,��)@1�D#1�!6�zBPњ�9���0mV���9iı��1{:{���B�����Iٹ{�k�L�/|*&��=P�C��8��g�|�)��1��c68'�p��s�����g���3`�����b`?`��0�9�,{V��y=I���مD�yqo����tp���կ�#����~�~G����)-?�Ž�^޵F�x��\j �B�^1�a�����G��R�Щ�:���N��F����?h�v4n�u�k.�6`E�Ʉ.�ѝ�j����|GN��,X�VD�`#�DՇ?�����w��xӛ����̈́�/�N�`;J�#64��f�Xf��惫⸰��=P��l����D���a�;=\6�e2ˍ�����I,��}D��+�(�yh�IbZ��Vz/��1�ZR�^�C�E��XQ��h>��r��C��,P��J��*(N�p�<��,p*�f��?Wț�ea�8yJ�M����� �`��s�;��|��dqds��� ��1���i��� ���F>�=L�����[z>Jέ��TPիr���A�,�$k0N�Cr�5����ú�0/b����"	,�=91e�	���U���I���p�$q�t�I4�ߍ���X�e�2 ��dŊ���Й78ق���k?��w1|8'��ߩ�����r|�()X��_h�j�Э���q+�D���q|��6�����0�ޜ�W����(`}��l��Ij^+Xb-Y7�0�C\�)���{�� �,H��_=���{�Ռ�3gB��������[�:����\�0�G|v\���p�?>>C�|���S�g7/��J��珠��:#E�%�ߢՇ�b-�o �d2j,�l����&��8�,e�dB��ϲ���{b#h��u��ۨ���?V	�^d}1�0m�� �;Xh�]�X�hcc="��x�ܳ��f�=��C�@�x�Y� a�pQ�R���̑l~q/��(nf��Ru�h?��j�q�)���KH��Й�}V���%��;@ZY�R7��������˾��i��L濓�ϴ9tJ&�vt a������)<�P�<5�����o?gp`�#Wt��Xx�� �\g&��D0֜����3	�3p�����Hl�ÿ*?�M���8����l:cs��17��ʦ�4�e
�,��!�Ű�M|���,�<�߮/�p�=��a�{°�	�<�.����u��3���	�`��&��ǉ\�9|�;�� TuA�Z]zR���w��m�W�@�$��� 7��o�/}�K�w�ð���c0��_���>��ǥ�ǩ=�}�C��
a[`�ִ�o�qӷ��~��k4b���t�7�ik×ʹ�?�8兿�C�0s2�sq������`��ۿ�[��9����p��C�dl�H��!������g{L�F�
lME���j�z�=~�G��>L�'w�3LO���A�������� �+fr�
�f����9�F��D�I�8����6��)0��1<?��G��虑	����d����(L�g}�b�q���sz;�<��6�����Cs���������W���y��<������V$�O�q�8�HY�|O�3 Ny��A}<�`6������b?�O4F3���P���ΰ6B�D�l5���������`��,n��(\�h�}�͖}̤S��1�n�3n<s^�1��;!���Oo��'�s{�c��ii`�u����`}m��Ux'#r�ۢ�+��)�g.|���'�����M�4��h	�0�w��k�w�l��~� 
��
^
@=�io��s`���"�t��|@{�,��Ѭ����_���?}���Ж�-�F�	|�ٺjSP�{|�%ףUT(�ݻ�����B�R=�P����B|�,��9}�d��s�܍ފO[܌��B��z����MFG�J'��Dn�|�x^=(V�2\f?��̦������|�����x�,��I�XC�b~�c6�?9JGR�T+�����������r����>�oQ��lI�l�7\�1L��I~ ���Jȟ�E YR+!�$� �)�1`\0`\�1��]�,ٖUn�w���g��9����;�;��+m��\͜9�-��gW5�?���U+���bZfO�*`A�Ey����.1�l����[)��a�;�l�5�GaY���H(���cQ��p<�-���k��7����Y��{�ޅǰ�����"�{��P�4�y{^[�w�1~�����W� Vڣ�#�}c�+m���?��UuN�W��ZE*e�|Qq�^�-�w��m
c̊;l �����+�u'j����2y��؊S��Y�ąN�*�����8
��Mt?!c��D*d%�ez`�<m��1X� e��8�}[������0Xm��%K�m�p�Z���,��D�sT�����sl�$���.F�<�
���3�56Z��(bKgRzL�Z� ���#�(1p����JX�F�A!Bs��.P�Z�� � ����Fh�ز�N�b�(qL�R�1�B���9f%lR�v����G��9�t�b,��7���x�	���8�}.��sj���ϙ3[Fǆ��zp���A�]~��q��ߢ|�VK��!�дg�A�WD۱�0Y���}�\v��N���Z.)�b	Mݻ
�Ig����uN  �1 @�l��
^�fc!��Z��GX�YL��Iu�����&��N�Q4�U`0��Lm��u,d��dT 2A�q`�)Y�KfNm�V���"��Mgb�:��Η��,��d��r�S��N�	��1��2��Z"���ñ}�5�Ԃ9~�'��ٓ�<�!S�q*
y
��5Pج¦���R����� ����պyO[0�}��h�A�ь� pOj��5HAa�/�OXw���7�Y�
>��,=�9�u.���Y��sf͒׾�5���\���^a���S~6��4I�Ƅ`�g��`yL֟z���Ȭ�3�f������=�ec1\��c����9�Md�6ky���._���b$E��� �a���B�Z�&��D�$�؁��K����d5C
4ݘn��Y'c�8�#0�!5yj�d�8?z�W)Y�O��M�sw��59���ٳba���иy��[�%
�;�.BQg�g��92�����b�3\PL ��X`�cQ� r� b�>�bT���xˠ^-�������G�f"K�L������L�������a��D���&������cl�P"�Nz_�����t����]�O�tQ9!��U���_�����%�8��ݷ�٧䷿�[��t캻���h�)9��c��7��u��k~$/�� �@z��ml�i��C	�z�8y̓/<_�͟-��N����~%[�>+%'�!e+���9&O<&3,ǝx�t��ҎPhG�~lR�?��]�SN9E���_�m�K퉌����$���"2C0	t.BĶ\�ϟ�-�;p΁e4ٽS_�j�\v�eu�t&��Ʉ�&��ǀ fs�A-���.���Q�̟Z�O~z�jRV3�1�
�L�-'ў�`iDs%�0 ��o�a��Dc�p�b}��K���.���C(�X4����C��U���M
e��s�9G�=(ȒZ?^�=p��z��x���S�Źѥ�!a�R8[��>>��kY��f�{B;�3�<ӯ�Tz�rD`3��%q�/c�A��ޤq.4�w���O��|`\<Hm ~���uD�� @;̕+�;!^t��O6��<������(� �z��k�rB����M���;������B��`��� ��YS�  �A�-���\9�%R���}���e��s�;����-�����'w�u�l~�Ey�;߫Z��@�>9�(�t�^{��7����_�z�h�� ��_�<�7�abc�'�	'�0�1�Uc5i=4<S�����8���<�+
�]n�yO��غ	B�q�ʬ���jo��0�?���4��P�h�y�\U�����f�02+�0&`Rt���E{>�#�9s��r��hL���)v�^�����}�m��*��i|=���cM���E;�ItS]�c>)�gŊq۴�������Bj7#��&�׮�S�y��C��82ִ�]?6 ͽO��Z����ZQ{��1f����G�޾��o�J	��P��k�S �,�?z�<��S��9�;��~��<������ʍwEN[�T���=�|y���Um�|L{�6���is���渍}�G�s��;n�#W-��;�ir�ed�_��7�G�B�� �<ޠR��6���>L:�p`� &�@7h�hm���7�u ��6֯����t�n�6H���b�H�9��[_2!0o��Q���vM�ic�Wۀ4�),,tv�����b_./]td�60=Q6�2dtn��|]O���0%�źk+_p>WPE��@ 
��1j���0F��gLJ��͞�-3�5�y�:����S+�A�ҹ���x�Y2ѵ�?�k�
,�Mco�8�vp�úB������WW0�� ���|򓟔[n�E;�q��~a=�=��?%�g��Z(7=	�(�+ȩ�Y����W;
._v�
�#�X#����[;�)W�N{��,ϟ�L��×����twed�K/ʑ+�Ȍޜ̘�U(]��LAd�Z��c�ve��21��܅	�f4�|���Lr��.��b5��XsP+AýMt=�O�m8������l���7HR�M4�z
�����Z��q]��O����y-�O�I��P�4ux�
f��x2Qjy4�q��lf��d��k``� ��x-��6�)�`��ٜf8"�}#�$÷)�d�xv4Ɂ&��r���B�)����^���Q�̙׎!���ϛ�}p�����Mg���|�l�5쫽�?x~�g� pK�.U��������Ö���B�p(��7��`�6�>"�g�d���2w�wÏ�X�hA�����-ȝ��[/\!�3g����e�aK���Ti�3�f�����F��;G%l��-۶=�-HA;F�v�;I���[yL�|�8�S�`�Ϛ�AƑꈺ
�����_�1����Њ��翐����̙77�Y??Lln��I4��t�������y�|��Ǖ�=&���s�E���q`�b����:'s�)�d��]�
�����X��6��f3ڋᩧ���$�;�L��ܺZ@����70(���������3 ��
w�r���)�C!±��êD��fy��6&���঺t�z���?�-/k�P3��q��d����a�ARY�.*úRk���M�m��b>���*��C��MoR�/�� ı  ��s���^{񅗜U��?�(�g���NȎ��q�"�q�Y��ky����.�M�����_|�y�Vp����h�3�Qbb�v�ʦs��Ckԁ��lJ��ɡ��c�5�ӒqǏ�n���Q�ƄM�F�^2w6��d��M�l�9��=a�a<�,��5*���V����O�qܬ`�}um:� �^��8��Ա���}c������cj���6va��Y"w,	0�fy�,X��F�<��gצe����%ƿ'"��®++���I����"�f�q��ʰnЫ�3���|�󟏳�p����ަ�~�/��8]'N��#w!Z6VkN�G6W&���J��`�qp��)�t2���5�6':b<��O��B
d�8�ȫ^v�
��g^�Їv��wҵK���ag��iSK��;�ͬ�X��p饗j�j��@0��{�y�7d�gf�X_��$n4�dL����J܂�%6�f7>c��L���[�i}��\N �1�c5P�l=)sh���8�3�+��
U��-�i�67����%%�k����c��4c�v�9�|>S2Pm����#�wؾ���xnd���_��j��v���������g?��c|i�0#��B����3*�rF{���ު��yi�Q�@]�iY��-�Ҡ����S"kHR�0Г������x���	�_��	�/=��=g�̞��i�nӧ
jrժ6 ��K���\�Grd�5�ό�{�G}��}�k��;�6rva~�+_����7�f�Y�n�6���Zs���u�-cO.�F�d5�fZ0�ϑ<�-@%���Lx�d�Q+4��B�g5|^�~�8s�h�Xo2��˞�ײ��^׎�i(�~3�k����K�}����J���L�eb���e@7yO��ܛ�k��`V���뿎�'�� Ա�Y���cb�
�×.��b5-�l |"B5��I�`����󥧷�E�>�E�B��[+��q���?&o��5_������3ϐ�;v9F}���}��9)�#�fuG�+9YԻ��Ԟ�.+V���-$9Z5R+����P� r�!>����>�1�җ��ھ�ٸ� h�l�7�'%�o�_��%��̈́�ua�sY��M��Y��t3q��2jF�1w���|�y�6Va��V�?��y�ɿ��������
�f�׎5��H��9��[?=�����co�CA`c1��j���]�E��MaGK ��9���{����p�����@	��dՑ�ep�%���B�L�vVB��U�Y9��3���k6�G�@�>�X���$޳�0L��P�����\Z�{��.7��{�L5ǰ��966$4fϤ��v��r��r9�����0�M�6�@N�h,��.�*`��?���p̒a�������,m'�!��Z�e ����2U�:HZ�>�L�j��Ѫ�Ԉ�l�E���&�߼n+���&yV��3
C+x,��cb�Jj�,���P�ot�V,��{.�Z�1Ѽ�m���B���(vC��;3߬0~�ޠAw�&p,���:J��,;���T�Y�R)�M�1�h2�ͻs�e�;�s�tǮRK ���[�QQ�k��:o�WUZ��r��r�mw�+/8_F�Z�d���"�������c
]r�I���^"s�-t����wOp���_���wj��~�� @̶m�����l}���bd���w�/�9��i�$����ؤ�8Y�����h�[ �%��O���ǤO�5b����`�2+k�7Ҿ[y������3��cac��ڠ�T�2�F�9?�ț�[]TlƘe�������v-���������KZ�M�EV,y$s�uI%�{��塇�SO^'��,9��N����]���������b�r�y���k��r1����]�=*]��b�Dn����?�?I~� �'��?��P��c�s_����\�������ŭn�f���9��8�U��� ����=�,���0�9|���*�׮Q낛�n �q�O"^�D���Í�{�I�}���=�s翭��U��H�p�m�)���p{��>R��粩�I����
~N렙�k�u[��<&7�s�T�Ɉ�g�xr�W���Z���fa �?��?W�>g��f�� H��;{��\�J
�9��3�UGɖ�7��� %��L֬^�, �SR9�%��#���?�ŝ5.��s��V��=�oF~��9L��\u��w�Z��	��9G�Ξ[߬nB�ق���u�}/�������?��?>G�=��ƍ��͛b�.d���.Y읤o�L���`l�2�F ɸ,�� �����>P#�ОR��Z�7I�����ͮm�C��7���jF��1�&��~��o����a�k�m��k� �}?p�Dw�2��ـ�����A��
O�������7�M?��gH�[����I'�.���xP�]#x�P��n����:+�?��� ���S|�����^�.`g#0s�q�)�6�}L$.��6l�GyL�=�0���l,�w��ݺP�@��8��?��'�.�={v�;5�v��� �8#i�X�8��QV�>D��`%�ka��}ٲe��|�f=��E]$?���!�ҽ����{?��b;�q��b�
�'2��/bk
(N���=���Nhx��g*�B�z�N@���u�W� S�7C�vI��}� ���u� (��[�@ ��>@j 4���|�Wj��Ƣ @�> �z�ߨ��XP� Y'���
�/Ns���Q0j �vb�:�S�a�#U�C��Z�@�E��x�`�Ŷ��a�Ê��������C? �;aR�g�2�*j�V��R�r�_����ө��N�N���G0�Aq�"Xa���&
�
�Dj*�7Z�����& x!ЋB.��~�a�馛tB�����f! �:�����Ad�eQH�F������Ƈ��Ob�������ܢf�+����˿T�
�u���� �l����3}'����ξ�}o��4SWÈ��aӞ�7���<`pA, �xV2ٌ]@�����t2Ku@+[}���h�$����=����;��&�M[#=��"3�=D��`%��2�M��1����������` ,	��{M�E+�?���� �֮�����[��gS�q�FA:OL�g��|�8�!���Zq���.��-�3+�S6�[ڝe�������XT>@�"�EĎJ6ۢĸ�f��%����{��E~���v��!���p�0����}�s d3�\�f��dVF*^ڗ��BOlex�>�k����PZٞm�g3�OGn'���R� oZ{�z�|��K�4���E��v���_�O�ӊ� ��XLHE��׾��* �o���ЮۅZ?�6����l6������=n�OX��`05||��O�~��/����f��|�+V|L�1`��
�y�@N�{��LZ����'���D�i�	���g�M�����]��N@*=��"�Whְ�̜Z�L>�����҂�}���"J���4PJ�$FK�f~�h��)��ŋ��� �������E�<���5�O�8hNcކ��ֻ�Ѻk��`������ҩП����/�l���m	2��=��f�Y�E�3�#�^����7[�kB�q��>��<]�A��{K=B��/��h�	�+�@�J=��~�z*�׺�ƶRZ�D�02��@<V��oP� 0bҷ�ܡ�$ѯ�ģ�3���(��^s��=C�;�X��e�M|*���y�X���cŇ���@d�X��Np�=�j��e�,�T}+?x>�r����z�����β��J���촞,Vp0E��^)'L��3��� ���ZM��N� �k�]�ijn��1����� ���[�)����U�xR���@�琡ں�d�� (�$Pf�AV�K֊���bƎu��,�m��?����[z��]��]�"~�N��sLg�S�����L��aJ�����[�!�hzІES�g	�,w��ò� N��G�x�z�"��Mz�p��DGc�^K��s�0��շ�yj�48'�o�vl�
ٜf̔��fh�K�k��cJ�RHd��E�ð���;GB'�*��ҹ,L7񚿿�={G+Č�`�Kѽ�:�e�J9�-��0�}G�����/�K�_���71H��t+�Aºd&W���@!�%P���s����O�Ly<{e`�����R3EN[�"#d�5~>�,j�_���ղ��T�h%���󟴁�����5�)*W�:I�5`/GЭ�jݯO���:�m��V�"s�����M�DR����A����YRp�*�����O#�F�;����>;%i����;�̌��B�t���<t�8�T�u�A�,��|���쳲t�ar�y��9�,����NP k
̿
�B�1�ZQ��[u���-U�W���H:�J_��|Ӎ
ّΠ�O&������q½w�*�8>��F�,5��}E�_0[Z�!�M��(`�x�����T�|�[8��dd-�F�t+�L ���5x�*nQ�O�[�,�EJh���i��C	�b$@���ה�����3#n��H��V5���v�I?i^'K��6ɓ�k~x�Ө�ҋ����n0f��i/�]�E�Z��eo�_J��ݲ`�|��;�i@�R-"���4�XK2�Ǚ��;�4�Tg������E(�� ~��3�����	*���䶕���fc�nӹ�̘�#��,�o��Kp;���@�FF��B��2P$0~:P\=�p���&�L L�%���SH4�R?�J�e���GX�z���zu�R�F��z�(�<nw�Z��k�!Ϳ!�}zٰ�1�rMq�1��C�n�u�.����(���}n���wO]���mTQLַc�{Β�YrQ�?�}�i��%g�h�Ϩti�W�� ��,�h��~{�/��Iw���Ԫ���^ɧ�B�He~xǂk���!��.�9&0�"NVkS����g�?W-�� ��T:$�ZY��9uE�
y	�Z��Q�����"�XM�ʽ8U���Gx�LCf=�Ex%fՁ^����
�6k���Z]�&C�X��w�8X�*��4Ѱ��������5p��A�=4|,("+
����n��w�1�Ë��M�����	[���b2�}���G�9F̐l�G��Uefź�5W��xn��3��*B�^Vj�蕙s�h���`���%�<:be�7���9���gܳ�z�%ǐSmdD��i���ԱgYcN<S�FS���	�J�397�9't2��S�b���|�ΠӚc��D���0�FOk���`�׶4���E~�Sr�'�1��؈,�?_+���fb\��B�W����6�ӰKQK�\1�������>�h��[�MY�l(�)��ŗ�RN?�tQ=0J���>�9�u���jr{ٮD�dU��Pۣ���Į5.�ae����$К��������1�*�����o4����vz���hmX�8m>���T��y��s�Nh�Kge�1�.�}%�I&�չ��v	�4CrZߝ���
��sK�{�.'�rRvB�\)�X��!˖.�MO?�kb;4I�4����9�:P�%d�̘�#�'.�Ŝ�3ئ�:5�3β>��3��sϓ�n]A1�
�`~u��ZIL�������}M{���3hJ�ޞ�����sΕ׿�5Z�U.�jZ$�%�"r!k� Z��|��_��6m�tO[���i�j���+9F��c����qV����U  �"�;E��ct%�}���p#�qi�PkN�h��H���tI՜�VH���G�2V��ʘT���v�;�0�B��˘ȔR=5[��-Q�eU�⳺$����L*�Wh�1��~֢� 1,�c�����u2 69gS�|�Q��ýv �Dֿ�72Yy��ީ�������ݏ������w) ��UGʯ�k��m��|��.���D_L{���(f��)��"W��M�Q:��M�T�n���"}�}�`��Ys��Xy��dg�q����ۿ�[\-�I�$����?��?��~���'�&�ැ�>L՛����3L�Q����n仫pH��X�� ���{ѣM�8�B������$,�J�����R�8�;�>K�J-3&Eg%Hۚ��}G_�'�jydB��H�+�Vk("s>@�T�9�WM��+O�������5P��n�U{y�`2c��݊{���P�t��u��l�e�{��J{'��I��� ��Ś�~���mJ�e K�{�ʕ-��P�9�����K��a�ڬ?޳���1�������6Y�z� ]�/tV�}�<�ݼ0.,�#�X��u؍UY���Μ��f�k�<2�n�3��ɾ��x��*K�,��^y�t�s2sV�lټQ~�>y����o��Du��'�g��Qǜ �ן����e�]����s�9��կ�a�� ~�t��o�]���oi�7��Y"֠��h�M�{J��:t�F�J��8���0�i��U�V�-�·��L@�&�]x���>�.�2��Z �4�`Yw���G�1��%���R��ߖi��Z����tYw�M��.ٚ3�L�%�J>�M�`�<S-z&]BG��Y+�b�St"���H�<@� �
{�9�����p��_�=�0 �/��r9�5Z̈ڢMO>��Z��9�:�v�nY�r��~�ٲ�5�,��;Y1�  l��Tb�Ӟ�7#g89�c�`h����Ҷg���[��#����h��Ӣ�����V����}�yH=��3�_ߩ�`,
hӐ�-^"7�|�B�b°@������=��3yV�/j+,m�7�Oj&)��\��(�pZc>�6t5#���K���s�������ˏW&���VI;��7橥*�ʨ� ����^��� ��J�$�6��d۞��m�62(��j{�&�M�&���70��ɸ�M���?�LP��ReS[=K8�N=C������rꩧꞇ���/��b�����=�ZE�ݬ8��ի���O�տ�rܼ�Qyⱇ����+�?,�-c�J�������ΖSן�	
�7>����r��^'t!�)��g�M*|�Y��*U��a��淿��yY�l������^ �<�B�ᑊ�x��r�jY�x�Jx4kA��>K,��[��Yg����������?_@<�І����tM��{*�aG�Qq��|v�P���@Z�5rbld؍u��AT�&��K�?��?A2�j�pM�R�Z��u��b����1�q�5W��ـ!u��+�Ȃ'2���2:��0%�{��G�s[�oߩ�C�c�ȯ�JH�H���%3��;:�&�e1ЦA����*~��R;�1J�C|�d��?^>��O��c���Au����~m����^}�,�x�*�]��2&�f܊*h��wUah���䦛n��K����T�@�`~[p���nA�?'���eK5�6�Ч�yR֟r��.[�̲�8������;�\�J���>���;��|�n:�k�qD��"��w���՗�n��F] X�X�����$�)n{N�l"��tE0�6N �̘׿�m��RM�-��*�28�]
��#�$��|4�ew*]S=� R1��B�3��0��V��!H��ޅ�S=}͇w�x! �P�RtLi�c#���ޤ$���j�I'��4A���?'�4�� �P����:��q~��~}>�ʗu[��x����b�Y1�2|@r���2]tP����	���к�u�E�{� ����/|�ʨ�	H���ʕ��yxý�d�Y�h�����;.М�+����s,�����j�W_�Z=Ǌ+���v��V�m�3�fD�����ӧ����s2:��&bT*U=e�\q&fyX���� }+����I��,6Ӯ]�T@@; ��{��^��0�&:����l�@�|e�@�t&u��$Ԕk1��~���'^>�rԴQN�<&)7���ՃYb��`��s�"��? ���PqO�ӵH��"�Зz`�0���T �� i�C��F.�0�Ɉ��9�8K4ɉ����,�KNͺZ?��.i��F)d� �8X�\�{ҵ���<7����ۥd�&�O���x(rK�.�7���կ~5{Z`���Ν?~�ȥ��m��='�4�n��lA^�a@�c:�1}��}�=���/����W;�0,���k�Z Ӟ�������g�%cVq�3jv��	(9T�l�riDjUg�� �3�j-@*��ɬ��^��T쟋��O�S�����MDs��K����[9t}�"���BA�cHtu��m"�����h���͂^
�ﯦ�W��UV<� 5����%��DA�v����Dh��T�sBp�v�g�����^@���MnR[	�,��-n<�%�y��$��[�&�̶K�G�;��y߼w
�����a,��If�gc}���+�}�ϡн�oTW.��ڵk����C'�w�Ճs ����~��R��}NX��Kh�@JQu5�ᾃ5��R��c��S��i���5sa.1����TN�xs���������� �����G�)Mgh�0����oD���h��Hjm�ק/�M�1�8��h?��f��>7_ǄC���Hۍr�c5���5��w�g.�CuL����!��(����
����gS#��S�o���#_��Pg)�4�S��8rt�(�ã
+h�M�L-�W�g���p5�����M��mj��NQ����Z6+Ǧ�RC��kƽ�p��a�C�>�ǴK6k�����L���%��O��
=���NS����}M� ��e�ݧf���W�������og+I�si�	�2:6,3zg9!��1Z��JM� O{�N���4��]2:R��+��KfΆy��4�R)#]��NW4ҷ��Ȁ/RM��/���1�!��W�*2!R:i���X�h�UW�}�&�d�%�.�OM�����2���̛�)դ�������	c�"恳��+ձ��s"�240���,p� ��F-�� �vL����W��uB�-���5�SH`��J��[T�@� X.元fi�����r26<�n������QAd���t��y�Mx0Ƥ4VԂ!
u��y���� ����|���V��H �:�<���$�BbO	���^�����تZ���x+��o�E�������[������;]W�����E�:�(�\a�޿��䆛n��R�6��4Ȏ];=�������e��Ŏo8K��B�L�o�ҘS��&�/�X�ם�>��%�Ok��j>{B��BӞ����cOl��O<N�֟z����K��]n8!���M�O�����)�y�n9��T���7���>�nL2���ju��
>Z�數Mls�4��B0��dұ�b��N�F�r�i,��1~�؛׮�;7�_�j3��+��(4m�<���������x�1�Z��,��9�|V�n�T��L!�'��Ouų(J(�Jj�D�%��1�����J��r���u�:DQi�Ϟ>|*rxG �>�|��?u���آ��B7���;S�=�x)�������~�2k�B�(��E�9�,��v�ˮ�a9��ӥ��[�d[�<-�7=%��yiFmߠi�bM��0�P�q������Wʖ�7��%-ꁦ72:��9�[4K�=cr����J\,��^zI6m��4�L���ze���C�c �yx�[���e��D�����[<���F͛+����is�7	�-��)t�E널�H�<���x���b���{��k��KP� �Xq�1Y'ra�Z�g'�Tݴ �\r��C.���X4FS��f,�mړw`Uſ����ܠL��-tfKe|��������b
^
�hjd��<�%Ō=ya@!���lJC��'?����}�,=l�<�н���!w��S��d��T�Ȃ�K�R�ʪU���/W�cht@�{�Y����'�i���������=�������'+^�����A��'?���~�+SJer�x���կ�E��Љ�tG�|�4�p�򗿬���1����?�o8G3��

ݲn�:y�Wz�(���3����w�� ��K;w�=�/�n�VՔ���)�zqc��-�1�7`�1e��%U ���6�H�1��z���l�dr�,��F�v�m�]�WoF{�jm�"z[�YhX5�a�k�E���;����d���3&�̝׿��qj7>g2�7��͚��{�Bb�ƍHϟ��.9��u�םr�-�r
�f�UK�\�]
/���s�=�Y�0Y3���Ɇh�QOWs�"���_�d���85nH��{�1NS^�����i�ٴy�j�k�>F�S�1{�cZN#t��-��"w�u�8�%,x��(?\<G}��@�lذA#�H�1V1��%����u�a�d8Y63�L��E����X^1���%$������w&�3�Vא
M=�ˠV���/�Ɯ��%��,��ze�PU������vR)�j�=R^�=�ŷ���yki���K p�iphX7�:��(7]�t&j���U�}�L?��u�?2�Ps��B���ه�d��{�ys溭�-��~��Y}�<�Ѓ�e���e4&�~�z'4f��pEQ�~�Q���~���.�ixƔ�M�;5i�D��	#��������G����n�3w�6MX�t��x���#%�Q��M7��Y���?��?V�����r饗*x2���
�Bї�a����k��ry>�b�����#��p�t��h���6�{ob%��묍�'}�04l�!��2&��(/>����%ya��̎T�U�3�xr���'��3�>�<';�������0S��rJJ��t���������MU*v/�C�&Y�$f ����Q�����5�X �:R������D�R��P�|���hm��×鱳fg�.��pX[8N��s�	���Oʏ�cy��-*l�u�����R=	�06R��z�t}�Qg;M��x≲b�2͂A:&�VKI�1�ǞxLn��V7)��0Y���DÒx�k^����|��؝��я~����.�H���!@��Ru���j�2�L./�<��|��߈����,��b)����3d=�:X5"NۥޞY280"w��^M�����ל�)���$�	��������f����K*�U��x
�?��<�V���w� + Up�A��|Je:�#a��Y6�-�h��m.c���R�h� w��m��;��"�}�yp��0�];�� �p���9��p���(bo�xޝ�~��/�����V�i�3�s���B��]�9�����a�͘5S-X(���v3�]��eǎ��s�7��n�219�D�Ϣ�|`��|,X��H�p�$�7p=Y�f��C�=��(\��	��)bQD��!M�+��^�i�t̠���z6ױ`����Yݕ�\
n����K*'�3��҇�/�dj2�/�
|�.oqQw�s�V�*�=�1�uTS
5S*Pl��gZ-y����>�O~��'��Q�뭷j���ɟ�7����"o�;�Lxf�32tː
�U�V�+�T�`�=�͛6�s��
��JeU��+|a_s~�������QGZ�x�	>$F�ˣ����;�駟�A=)����Ro���(s{Y�?�����%D�V���3�tG�ԑ�j:b����ݡ��s���q4{:=��u*�����4+Q�^��, �U!��u�⎫��X�`�)�RZ���L{��)���x�P-B_��Zw\{a�{\CP$�V�����i�v2-��
�\��tF`3n�v�&.�)�դ[ (��<?�W,�u�r�9x1�����~��T�����;��P�
�7�7
���}H���'u�m�7!]����e�6 ;�v(N���(�5֨�)�u��Ti�R�
��ct���2�[��3|b�KVPE���.0,>�>�я*C�������MM?�zDqd�"��Ͷ��m�����	���)��5�`�&�mj����}��
��_�����>���e�M@���C1W��+��̰V����;0+2D
������(�m�ʒhU�ձ�x�,f����$i2&N�TiV��Q����;�
|�����a��YP������K����BRp�"	�Z�/x��ʑ���u���ǫZ���p�=�oV����2e���#�1�1'��X���7n� �,lD,@��p��#$�+H�0գ��(��[�����ׯ��E0��[�'�֩E�X~c� Ўc�k��{*J�4g���Ƨ��Z�lJV�-?��#d��B������g��WŦ��*�����ݽ*[�`tP|��`��[�S3�ռ���4{@TX�v�=5��A�'�GsX���D� �{��+��)�Uů皏B�.���f#�i���u��g�惻�o<%M�o~���S߱���ޠ��WH�[|�����ˊT����R��~���?92a�����7��.�`7��CVӷ���$Qx�+ΕE��-*�?RG�"��K��G,j͚5��!��$ԠS�:g�&���I'�$K�,��<�ξ]z�]���F�3�=n��A������(�!g����y����{$v����kt�ӕf�(���\�!�P�nӑ���h؉�9�s2���qI~�1d�5TZ)�̮`�O�'h��8���K�����e�Ų�[c��/S&���b��[^����Jf��9\���1�w��}}����x���'1��Jd��] M����?�~Z����&�?iER��4U� ��?��UK%�&�'R}� �糀�����8���?1q��j9��3�x��`m�r����JVp�E�s" ���~V <|��u?P�������O����_��3И��5�-�	9��g���.����C��lAl���0�B,\ &���R��o�y��q�Zf�� ������1ל|��˞�:$���#�v�
���h��&/���od�=���2�aЗ!�HZ�E� ��v�*כ�[�xOt�C�h-
4SɁ��"d��פ�<Y���q�����cQG��e���n�p�?;��x�y�6���.� S�����/L�s&�SS�i�������:9�c�o���8��͟�b !(f���\b}pS��	;aj7�ĭ#Y�x���,�i#��=�8k���� f<@�bQ'��*���@{�>�V��z������RKK��o�
١�B����z\�`��7x4�kLW�:�dĠT��ֱ��!�ݟ|�ɒ&c��;��,$4�k�'
��-Ȅr���wr�;����O� �j�������>�A��7�U2��2a��%5������.K� QK�o!�9�,*�ֱ{O�ERs��x#�_�f��e��߇l��g�}���ek�a܆i�w�駱�t�A�̔?x3  ��IDAT�^b��YٴL2
�yR�d�N:;��e��K�Rq�!2ie��t��h;tY�	�;����e��{A��B�;��ĽMal����g�F��_��EAPW�gQ�2�%��w��V|��hL{�?��'��(%w���b��	Q.U�HWf�T��er��q���S�b���Q۲B�fh�o��-)�*���2��)u�XF=�9��ŜC1�=dD��itD�*�cΧ5O	�^����5�r
!�J���w-ܝ�m����):^�Y��Vp6Ef�6��rkѻ$�Sѻ��lΤ��9�c�y�f���oM*(��1?2,e2)_���	+�5��;\3͘';e1œ~ ���uL���je|FQ��3
N��P-���F�* ����;����K����ɂ�L���+�?,]C��	���e�<V���A)� ��|�7�r|A*���3~�<�fn���$b~���Iiyu�7�@g��bE+q��2����hS�#�[m��G�Ķ����ٱ�������?������}t��� 
�f,)�fY�(�R��|j�A�B�C
̠�3kQF�z.�&��B���|�)�L��g�5{����m=L&?66o\\{FO�2�z���H�g��}���̦Y@6�+LE�ء�Z�z��`�z�S�����l�;d�螱��{�8��Ne��:���;�7v��9IE-3٨[w</P6�b���B9T�#V�/m[.M�ާ=�o��s���DE�:��A#�#��/>L����64]wf]��m?�mMlLl�v&�mۙ�v&�m��}�u��9g��]�]]���[g�֨ ���p�Z�+(i���Tߖȥ G�M�qdM��2�0'��^:x7-��R�af$eS�[���"*D_٢U����	�&uj9ad-Gv%N(BJ�J����
�ǎ��B�wh[��zZ'.u	3��c$��6:qd�l��&�%�#^��V�z��˚93�ٷ���g��Sq|ܥ	���ʦ�&�8Iz-/@<2��TG���<�߬[��X�j�jZ��U�������q~y�J4C��h��"]�j����R{rU�R��4ǣ����T��9��w�Ļ��<q�;�F^���.������LT�"� =����<4ƙ��+�����"�+1�>��T��$-�*��y�D5Vr�{�l�:�r�Ԋ±�Ey&�����1��d� u���b>�ѐ�N/�7AaU��R��o�tY1�7㻇X���pNcf�Ov>6��þ�p��wH�\��lI�`��I4�+�=�J��!p���s��ɰ�F��X8E�8�SԞ0o3Ĳ;(�w$�J�0�'�%v���
������ 9�:Lf�Wew���c)����p�"Ϟ�Ê����Xag�5&A�H�� !O=,��{�s�Лπ��.�ga#6�J�	���������-�%qH>Z���ϗ0_rP���R��٣�!��H�֛�P�E���7>�ic�����v��:w�:�I$W�kj�o�*w�[vq{��ͼDM(��ʗy(�S�}.�AO�?�p�����i2 X��MB`<���P9:�1o�}0h����6wp �4�\t]Q��@
&uUS:F��f�fD�*��y��Q�y�kSnq_�W$p�^�����Q��R����^�_�<q_�e�}�B	���N�o[3��!#b��V��.�e���	�Ȋ����~��e.�a$�j�\k�����l:�a�K�8���d�X��y��e���s���	$X��D����Y��S���p�?��B�i�)��F���Y�*
P`:RQh���e>��!�mN8�Ev��q��B6�~#����3�-F��������2�������ҟ� �R��U^��~�+�^?p�������濑B�����ݗ��o˂Y�Ws.a�J�b�Q�hT��'�]��M36�U��4C�'G���{wj��r��F���!`u����y��)U���>�a;����f#���UԚ�H6�뎛*S%�;ڼ<��3�Y<K�6��������C򬷟���d�=w͌�c����b��e��q�(_��1'@'>+�>�]�@���m2�ΜY���c*�x�z��T�S嘎���Me���Od��3ǔ���˭:h�l��1O�k%��S�:��쬧��SZ�ݾ�]?����S�ܽ�E�/�	�\4�M1��6_y���d�j���Ue1���ѐ��Z���,�j+b�4W��d�aɞ���D�����qAL\K��_@�q���s��Zn02��k�4�\�k��<6̵���[+&�$� �>���k�������� wf�:�V��>\�e���x�����*�;�M����F��g��K��;Lyk�����Fe+� 5iQ��.����4�������/1����Yj�4n*�����u*�֐��P�ɿ����w{�����ϒiF�7?=�h��.�bW:��Z��.�� ��U���ˬ1�x����Y���Ԣ
�W�ߤzB=Y�B�^_{��9|vڤ���%LuyU�e �-r��Jڷ���n����(�8��rk6��q�Aec�\�L���o�*��DP�m&O{y۹�o����8�3���Bi�H�~��P9�������/�*����3�%�#nR��ViӞ^0g�>D��,e�T�}�:�9�i,&y2��^�8x�d���4U�pQ�0��8a}�K��``������F[�2c�K�QW�n?���9�>�~?��nkw��-��������}_��}�8>�i���J�� +��L�=c
�+�X �kdw�4-�
ʘ��9I�b?F&�s��ל��本�">�IoL检�*Q�[|�ɖ����c����8�&,G��d�}wJ5
	;�#���q��t�� ��{�P��w�-a澜U�� ��@	���?z�˸KN�|�}���͜VK_�Q���?����ZE��~��}�6[���f�f��ߟ��U��0Wv���c��Ev��Q�	�YH�"�W&�W�B�xc�����RkV5�-��x���������z͊9[w�<����e�|Pi���R�<��q*�,p��*6�n������&��R��q�
�v�s�z�q��=�Uv��u��\�'�������i�H@7���I����ӱR�V�֋���q�$�+�Sw98H�t"�y���ݳ�|�@�ٴ�p�+Ŗ���P���u�m������Xzl���Jp�� ��B�m���=%����:��"������&k,4�}c��I KW���Y1�dx�O�ϓ��zM�>�zUn�Hv��/x�6�XE��S9�	O,�����PP"��i���(BZH�]l�n�"�Pnr0�i���b�o��$�Ѡ�j�Q���T��.��Ѵm�~�1>E��浱se�2^��$��w1��P�h2�Dt�oh6y��:ltL�3}P��<2����t�	�/��N�(��#x�bL�����Q��?0RI~U��?&[g�3A�� �M_F�I}7F���}a�A[m�/���ؠ�p��o�qD6-"'�_��t�_O�ze��sT�妅�t[ބ���؂v��~`��Pq�)�)��&�鄲�~�2-5ڐ�# ߫�D[��QH0�P��e~�Vy�I��C-�L��Lnk�6�a��s�7��}օX3o���b>UY�3}ف�u��ߟ�V� ްU{���@w���C�t��t^��w�*�gH���Y{iǑ0�\��~X��6�:��!�_6[�Օ3<'lߌ��>���'X�&Yy�4xOʕ�5�M�iDc���`���k�`�0qA	�7 ����I0@��w@@���'3��: �D��q6Ap��uX��R,�7qş� �N�����9{	#v$)�8���Z*��s� �������=�[�9�[yK/]���ZI����.D�܂K6�M3��,��r��G�X@lv]��.˹]f�S��T��,E�pQxོ͕K�m�'o�;7��\�1!2z_w�lN��������� ��&����v[�a����Ƀ��
�d��-J�����,�vUP�?�Av'���/-S0d�����l�2K�A�ړ���u�N�咕���N(����j]���O+"٧6�<�O�7��$ޝ���L���,^!=60��E�9��}���agM��%�O�4���b�ˁ�^b�H�{
P눻�#����v>iX3��#W�^3�_I��r���I�6�lc�����p��n�2��v�����4(i�n�d�N�ˢ�3ރ��+���Ӏ��řp.p���c3�]�b��]�5\'0���ۦ3�C.CS�k�[Ҋ(>{O�&1t�/��ȹ��f�{5'���Ϛ&h&���o�^[,.g�t4���?�cbm�P�%����X��'��ۧ�)z��
��7^��?�{�S?w�)LК�;Q:�3�z:,�13،J�toI�J���{7&1Y?���=�����%1�ޡ���V�p��Vè��M@����8��_����A�V�F)�ĸ�ު^�WՑ���*�.ܙ��h��c��|���DlJ�S}Π��ӊ����?m��,���T�&�%����������{�N�m���#_@Gc�ΙA%x�����6ɸ2���
�e�;���,��u�2庫���������~a�/x�IMyHvVb9�6�^��̨(\��O|�*���t'�l��U���=Y��?��P8g����^i?�o�Xy��3�"aZƟ;XGT-Z}����wy�f�o�侓-��Mq��lL0�R6d	�_�V��1$���i�c�OB�0a��� @b���2 ���i~*1���/�/I�M{�����O��_�y<?�xJ-DP�����qrb�G�ǂ�������:0��D6�:($�#���%X=�il	q��%���}U=�MG*/�~?�.�WQ���^w=��,��$*(?���.�����!Dq�*��NI�<��]�ǥ�T�8�7,F�i�����\�W��x^���+7{&����<�`��;@#��Ϯ�,h�/�s���K@��e���I�6U]E-�pj��a�58^$[-�3��.��e�$�������!ѫ�l�hO��91[=պ���\l�&@�u�2� %?�DX�s���bYow�����H��i��l�">V����B
�+0�[�GAKI8	�m�[�@�Q�̈́�X:Z�X#�O|B�@X�^���xwh��!M���E�q�QAsJo�e/гInv�{�������a�(Wi�5�>ig����}M:��=��b���W>�����Є�De����+TǇ�	t>;6�y��l9�F��v�6�������W$J^7K�W���`!r�Q}��%��ƶA�� �q[���� �A���M)�]�j�v���C�ڂ����ې�oS���bg7���C��|�خJ��}�h�=u?�.�E����Sr��T�ݸ*{�ݿ�%<:j�ܹ�o1i�y~5�Uq�d�D��kf���_�rAc�����śᅟT���I�}�a&|0e����?�6WN�t_Flr����1�y���?��(��f6�����7�[l�Gr#
��I+7� �Vk2~����L)��z�EG���x��W�Ӡ�~l ?�-ؕ(����Η����2"�2���ԩ��a�������(�Q�ffe�A1,�f��yj�a���5F�j=���^�ŃS�_����{|��ҎOj/ ���=�p�6�4ͫ�B�+ͬ�`��[q�MR�Z���S��gt}u�|X��2šT�W���#>� I�C�v�-�r��l'O��__q6V���N����Gw��1��x�����y���pP�Ӝ�鞐��ogiVģ�A`ZڻJ7�8��z^���H`�L74|������6E�P���GJ>DJ/\~6�]M|]`2P���q8T���lF}>�g�����6ZlFe��M�2�´�뿁�g��c�����Tڽ�z^�������s,�����|2��/
 >0�����mp��D��V���#4������ G��4�	�iC��Ԓ��tR�L������P�"�
S���ڷ�ڕ�&��<'�����{�c���t��ð.���Y2C��+r%̇�f�<�0/c����k����և���� E/-F&Pɫ�{:G�ifm�T]/����$_#��s�lBi�[��^���R�Eb$ZiF�(�#�TD�4x��F*�$�����p}��R��k�X���n��E�Gs�w҆�<���=��͚��;����e}Z���#̾�!4���)���	p<�v�0K&��\�M"G]Z���gf��?����%���7`h��.�P����m�ҵ�}v~���B�4�����Wg5���g��|6<�f_�=�i�;Ё�t`W8`}�� ����Y�۝���^f xsL�=��Y:��W�/�2햌nr�r�w���R�A�[���T�b6N�m�X>�6�.}|q�Εf��MPl�O�+�Y���R�oQ�l�U�.�H�����!8�'Fͼ"�EC����)@K֓��lY���q��H���;�^�r?+��/<տ	>Oěb ���i`�n @����`�!X�~�AFepB�04<7H���Fh�ܼ�iC���$�o��0*B`��oScU�<�K�*��8�B��Gi��'{�"��ί�+&B���V�`�j�����& Ͻi��*+�|���4e9��4a|�����������93D��;s�*-9Uܳ���$P�O�����*ίv���!��?V-:Dq�y�0�O�G�<@_>�nyo�X��D`;\L�9����xQۂ}�;T~��V@�(��4�ܰk�>��T)��1��?8kMi��Z8?A����y�D�!8�M푕�4����s�2��29�3L{>��q��3}z����8�-��L�Y=��@>�d�Eq=�BZA\\�s�;2�Zqbc�\�N�^ՃC�.�r�X��&\��ό��Q��@Eg�����DW���+!$1��P�O��9��ʟ���	����q7yi�u"���53Сz�����bs��U�:�sb,���˘\��W����!�{?5��c���Sc��y�:[>��4��Jg)�l��
�M�r���(�����&��b�@2�33�͠Q�Y���!��U����e/�\3@z[�5��4�+��MUnw/>��J�\IY�׃��z6E9<�F}ŭ���2K
��?
_��������#�lfE� #�k�^�7�&u�-�A�{5�{�ߞ�**��rI�$;=;�V�,��Z� F��/Pd@��<��6T����w��p� ���=���)�h�����'�3ٴNr�d��8=}�����Ue����?����k��t������G~�@�`;}a��){พ2ki.�R|[-,z�0�V���ex��/�2{��.D`�6��t�G�.��?ו����&$$�(2���M��l���O��2%<y~�,�s�I�i��;:d쫮C���[(�O9��KW����@�Ԛ�ݫy3nd\`��@�!V��>�XT~p�uá}sam���!*��F�� �B��2.���l��,��ȋ ��§[�7�~�YD���yj��Xn��Q��Z��ct
U׈��.�^S�g?/E����}%�	F��z������z�:���8�A7�Wg��2ݗ�E������d1z���T��(e4�#���\��a��쬧�<�~�Rٞ0e;6>�cO�8	����f ��:�y5X�R9��[ۜ?�%P�}�/�ҋ�	�Ve��]�t��!Xգ�[c�����k���!�th��c\m��	�EE�f��v��2G�R���5�1�π�vR
KJV�&2115K�T]Ϭ#I�������O��PRel1�&�On��N@c�ZcI�)���J�6��e���)��l��"�H�T�Q�V6�`ɼ&����A#��e6�!���<����Q�&;g��X��X�P*�+��˳"FOX�+��b�!L���Րd����(������p�G�.3�Uƌ�0T#f�/v�9�թ��0��|�����^+
���ud�]�,�)z�BOG���^��%y�=��'����i��u߅�*�:���1�i�ŝ�J�Tń����6 D���@�Y����&����+��(������� ����3�������L��DO�%+�½d�W�}R3;c�=2V�|��[���
�c�.�yf�B�BK-�X�А�s��s�+����MF��P����!NK�B������x�T�aӠ�Zbsݞ��:��e�%�;4�p_�v�0��ÍH�X�U���{�pa�jbi#_��	RԩybN����N�H�߼�y���"2��V���ui_�����k�X�]j8��w������F��~j{і����5��Ԅylze�S�{�P�P�9q��x�ۦ��Ɉ��ᶉ�ځhP����8\���j3g�K�c.G��h3�*W�a-W�&˦��/a-�Ȃqm~��CBZ��f�k�⦩E�5�A��10��h��&��!S��q|���t:5Lh�<8���P!�vxӻ��U]{�y�7����ЩyI��k+�&u��o�f݀��,���41�����;U����˴)9�q�1g���?��R��8a1C]����^?a�˶�� 6����WMDA؂�֟Ɲ�-�E"�W������������Ǿ�8�:��=���i�o���������|ʩ��'��,�vz�`s�(�J|lG)��џ�|u\�S��2����l������r���#.[�m9�<��%&(f���]�"#<R��o��X��1�ϥ8}�_'Mf�7��G�M�ƌ��j����*s�PR"3��	r��S��m���X����7��+���3SbV�	{ ��+
�fN��v���/�����/ΐ��Wl����SOP��_��|�)�ف���+t ��'m;�W����Ԕ'[Z���ο��h������)g�,Or�}}����~�]D?��+�fu�'���R������t���lን���< P��k"��i����jND�����$8oњ��ǐ��a��{r���r=�r�!��N���� ��Z��=�'�	��7À�x��vs&u,�Ѓ@��w����VʀS���N�)���V�h��d�C"�ĭ���m����y�7�@�N;��G����(�P�*Ćh�L��6�������;$����ʢ$�;�K�2g~�D�\�qUu�p|�*Q�]�5��8�	D����o�Yf?=gD_S�o�	΋ꮇؘ���O3&2Vi(��:+u$3��&�ځi������h���"vA'�}~,���sݏ�3�!��0����l���Eٌ����]&�9Xq�$f�]���h9`rM3�1��l6Ĉ� Pʔy����(PW[ n����u���m:6;f�q���7�0 ���B���F#�e_L#-����414.�sZ���0֙�`������VWd����kc��N�vӜ�x���
���z{Ðn�R�ya�qE%��r��q�}�,���L�j�"W<(�U��~�]�giդ4*�Wo<k�~��E+NР�g�>b�f,O������c� <�X���� į[�ѭ���1#~	ڞC��x&����{�M��	
&�d�|%�@'���^̞���"�!�|5 �	����V��y�z<�(kN�jj��p��>��`\ g�r��%�A ���y+nM�F���|.���{�I�L�-S�l�%z2a�d�f<��ǋ�<�QxY�	�%�'dn�K�-�P����֏j3�q�g�2ܿ��Y���1ط�Ƈ����#��ʻ���C:f�+ڶ�5+��C�H�ge��������}Vai���j�@ݤ�|Aw�q��K��Ҝ54&�ɣ�����)N5������{����4m�g��(`X�~r�H�H�\�����S��+P�4��ЉhM@��N�*&��o`��L�YB�����b���M5���"��׶�Ҝ��":�� u�'��[U`�_^��>_f�U���\�,V��������}Yu[
�g����a[?7��n������n�r#������F��ϣٮ[D-�O4�'j����9�^�E�O���:mwHeKB:�J�']#��e�	-yGK���I���yg�dm�9z�K'�x�����,<�t����1G�؆OE����2�:�Tj"99bDE�w������m�f��m˳���_m��1�1��Z���G<�@{kK�
.Ԩ�Eۼw�d�ctɾ��%pƃ�b�~Y�WTk��-c��
ED󰘆ou�2��]צ#*�QVK0����b-��*I1Ê	�r�+�i��1M�
9rU�hL8;�;٫�����c�^��ȴ��������a���(�}�FEiAE��h�3k�����faF���M7��Y����|�,B���)>�^�E�sU0�1_�	qrݴC�!�o��Z�2�%GRs]5/�X�]F�&>�����AX�M���g��P����[��:?3YLt���:vH{��R �C�b=%VQ��sa�^X�<U!��a�o�c������9��3��6w8v�"�Q(�\�B*�V6�\y:�ߗ�#M�o��4�>���ګ> �څf��� �����k��^����MW���p�N߸��n����A��Z#����8���ԨbFFn��mR�y�W�ǵGA� �}`���N�q�R*���L'5U,�ċW�L�ZiM��wծ#N�|���f��*�j8���ru���g�����ɚ��T>n�\��;u����q	��Ǆ[���_0FZm0��K���	���:EH�Y�G@�O����]=_���T���m�r2Z(zz�(E����>��ִ�o쨈�U�*���B ��[�lk��r4�-?��t��8�o��+'z�C_<�3�� ~@t����eveP��Ui؊#�;��B몀�^�-��Y7�:~<_G�E�*+�j4�G������s�~}r5�A� sq��z�������[��I�c�!�vhJ�����R�B�4��@G�c"�f.l�����jUbA��ݱM�����hz��ǧz�t�E��醧�N8p�!���ud��s4*�}"��b�Y<�6�S��`�����$C�(�JV�#�QD��e�TG=���W}P��tڼ�����&q���u��>�&��ڞ��dY+�|�)����&�D�_�4�L�Ԇ��9{��k��'D�	+ۼ��4����0�~��hd�u���g�{����xD�w���`j���0�(��~�޴y�Cˡ�ތ�#�w8B��!q�>X,ލ�Vz��������O�V�P���v����5�x�ٔo�rY ��&%d��X�qm/4#�PԤ[�����������K�~�V���a ��%��f��f�l�y���g��Σ��TR�gE�.�m��-�)���M�u�w��Ix�+�*��l�+�iSD>{=f�X�
/f���V����#���Ql�>���6��j0��5h��E�~��a�����z�W�����M�f{ݪ�JL�tqp+wK��]��觰�:m����2p�H1�q!s�3!9�����u�y�k�/��XZ,s_���|��Jʋ�k]5!�8�`�e�Ì����b:��~'��Nu����ʍ�ڻ�(D�
�8�x��܏�G����U��J�Fa	4j�i�`����1�L�f�P�Z�YOxĘ�B'�?���,��S�D2HR-�_���0�����a�F����jn;�r��~ʊ�Y?�Pފ��#�J�&����pe�� I8oo4MkRp�;�4��,��S���ͪ���l�����Ѭ\ ���Tc�H̦9+�R'շ7�����8���Ź��A����A�2(���F�\�;��!�4��ܯ�܋q�O�%VR�i&��!1D���~+��z�9���i���j9��_����V��0K�<�3[�9[����� L0���q�r(ڷ�m<t�φ5�=�!P��(gN�^*F����d�GN6ĺ演�Q����w˧�ޏ�j�Ӷ�Q���4�ph�L ��	��w��1����ݝ��"��.Y���$UL�R����O6߸@�=����X�˖F��@���R�!u��v�+� ��x2���(���g�͸ �qZ��P��8�	ru���-�#���~�#>��3�jC&2�@ӟGv�C��lV�w>����5UM,��+�4�M�`�h��R���4���..�I0f�?�,nT�ϖ�>4�[�<x?��}G�%U���0�D��0=馒����Y�4��t�lF������ ��k2R�Ԥ�^����GV�~���O�'�Ŗȁ{`������?=4�RzخAI����\ZCEj�ϔKϡ���_�sUX�$=�]�>;nfQoP���({��܀�l�H��՛�w���o�&��_�Aq�[�н�Iݟ��kxG����wi����F�B��KIh�o�S�Fo�����q�7xz[r�{k�˻N���@wN˂�+{q���Oui&��*ٸt#�LpŬ/���L�5���W��xبN;�W�n�'��*̗���֞�����1�*�ZnUt�h�ZӰ/ǳ
��/R� ������P$Ɋ���d�f��,K��Hj��Ll�rQp��:69������gi�c/̷�Z��K4*S�uוp	�땮qY�}kϛ���:���dD	l@g���#��E�fq��Tύq�s����KU'(���Q$��t�zws�"oh׉��F(V�MC��x��j����+Ȗ���5�j����?s����hu�,�0���=��\}=��d�
�c)>�&�����d�칤�]mҐxc^��V/tE��}t���aT�gn��~���kͪ��`����X����h��|��QGb�{9����E���cE�Z=�U�����Ø�C�C�e���K���k�0"6�d�}hʱ�}��5u��TǕ��G��\��A��K]��=��h�]�l�E�[_1+��Re�Z�ݢ�]ã�m=�]�,���
��]|l�coyiJl��	ǖ�1�VN+E����;�7$��٣#�&��`J�!bh�^���`�����IlW�0���W�3�ƺ/��q�b햢��ũ:<�MS�I��os���L����qFv��~���aDmlp:�Sۊ�pU�0���U���W�NC�d�t>I,�ě�����j��usi�O3a�1�j��gc�Z�Y�y�9c�U��mh�!�7 R�e��v��W*��<���滻J��\FrR���b/U�����*d]g��M�B(�K���L������s��'�(�A��&��=�����G��_ys���S��rW5�]+���e�J>��vI��.��MJ͒JM���F*R���[���f��+d,|Qee�B/��=kx�]���`Ѫ���9��uCX߅��k1���-y~�%k}�=�@�x�!p9�g��=��́���!��`�����'瓮�_�x^�o��@��'ұ;�u�D�oxS�rY�k�0%�g�^��>�h��=�#.U��_ay4�}��R��F?�J���}��rq�D3�BN�:���[��$���o�E�����&��d ���s�z.�7,"��������Ie�9��J2�fqLR��ņ�&�:�E��{���3ב�*���ĭJC/]��fd;��,J���\���
�5����{O�H�%>�O5���ҁA+�m�mB�8$�4�e�*}�j+�)����{��s����g�y���7��r=�z�S���pl�rϭy�z�#�׻F���[/�/f���R��m9[s-&�1��/R�%��l9�D���%
h��e۰#�u�kB��t�reM}[x5)q� '���sGӵo��R�n�|��"��)�{��;$Ӷq�m�c�Y_A���F������k��v���O�nxLg�m����"�3�*1�Z a:���I{�L��Y���kX�5���-�b	�	܃44�R�<R�׻�4؞�G_������#��͉�a�;̘���l4�ݩs$��kͮɾ�o\��� KR����v��3T8D�m꫏�Akc��TE�n�u�}�@Y?��}�� y��Z�4��c�)MG�ї:���=\�c��J��eV�� Q�	r�뢞��UʥOs��꿼���.Еo���z����t&���9/G!GJE���$�cfb�t㻗��b�(���Nɧ{�L�²��$ط2\{��	X���<�8��C��1 ����J Q�L7u�_�n�3 d���C���ݻ6�:��:���0����<�K�x9��7����w�jZTn��&�9踰a��0����ǋ�T1�����@|���8ːy�[M�Y����g:V8ݿ�f��F��[��r[�G���p��軨�y��˷����QP�ˆ���mu�3&Bf���o��d���0\A�΄V�@Ƨ�����Ӓ̋>Hg(h���Xg2�ix���}DO�4m�x%�̌H�����]-�?�Idր:NPTP�\����5�l��ѠC�YC�?:����~ޠ����u��y�y�8�$�;�+D�8����c�a�(I�h�c�;��r(Gcs@�ĵ]�+���%�`�'�>�#��4ٮ��G=��h�W��Ψ���~�~kW$	�q��x��.��� �m
Q;�V4}��,Ű�;��j�*�*��K�I�����������?�X<s��(�v����ʻ�sBA|���1��oY��}�'m۷2��f�V7�43��X�m������R��y�{�tbh>�CG/DvP�C�M#��O�at��dy�N<�ȋ� "}���L}�0�)f�� ),��0:��6C�Ҵ�N�!i����Q���d-�ؒ��x&~..]R-��/��e.����b�[�E&+�{;۾s?	I7���#P�ߡp��'�{��;�~,`x������6&Vpg�F�����\Ы|f��3W��؀��n�il��Aư��b� �j���f��k��92F��.v���ya�#I�g��m��_�*�����P�ߕ��a�^<�89"�A~*��J_��bf�Qҧ)[�i�V�+3*�z��*O���2�r��y��m�i�<,��%�྿7�Po�`�1(��O-S/�X��v{�M�]sC�zw5���Yt+7*Hb�㾤2�À�O~ZЃ����m�>%/�ZyZTw)k������K������j6��~�~>��b�@'��35��hGAB���ß�r�k� ����N�h_D�~m�g�"�$\��\�/�A�I=���\Da+���������Z�W��%�ʕ^:�I9����ȷ3eE��6�lRҹH�@16�L$�P��Gn�?�W���kh2A�^�g��$x^7!�&�������� B�LjA<��"R{^y�<��<N�U2�z�Ê����ɚ[���V�~:+��}|w�1���_ݻlߜ�XY�B�#A�,�1���'?�I4�S֝��3#���}�ヶ��k��ֹ�E! �T��?Th�'�/b�]�����R�*Vx��T��uXB0o~ ¦q�"5M�ɫ��os������%�(�Y����FU�����/��y�r��DѢ�J~ �t�{=�^��$�	��#�_�� ��E�ơ7����ҽ��#�EFn�ɸ	z:RU�oxx��X�?�06�oZ,4p��XY��~���	
�Ӈy9�%HkĄϑk�O���79� ������eK	��!Reo��a�'[l�]"��%��$�(�)A:�%����9qRl�{l^,��<r�-_v%�R3�J��2�╌'U�Oבb[�G���8�
���7+�fء68�ɅĠ#)�B��2L�6e�R��}�>Q��"�V��g1G�3I0f߶�qݱ�Cς�c�7VOS���ŬM����cy��Y����!B���ɀ�1�1�����v�����ro�Tۧ�����\�4�Ut���֣�g?��?�����\#�>�9� {���K?����s�A�����`�r��u��� h8U���)n�Y�N����R�]h�*��*�L�+�m}5���+�_��%��*u���E��9F���y��a����L.z�Yu|2fͮ�A��&D4�Z#�)�<"��䌦����'�&�A��xX����oӑ���I�FB���������5��|��0zw	t��7�N�m�{�仐Z0Z���h_����;��w��`�G��T8�O��������rZ����c"i!X�����Du~�he|�T��d�E�3\������eۏ�K⫻i�g_���ޅ|�c���mqY���Ѵ�>�*8�qX�ȠZ�f�|*Ԁ����O1��Э��O&��qᅬ!�^f8 �b���]����00�xՈz&S�HmXkU��~���w0>%qP�U8Q�.��[�*<ބN�v�Y0���xdg�����4��#L�kh��.�4����#^=Q��6�
9 ��o��L,�ߙ	k[ͳ�Z���l�CIK��]��=�zN�V3L��<# �6����/}!�(�QN�R�Gj�4ǟ��n@��w2��
�,cջM� �cRxB�ݫ�,R#)��W�m�����}bu��s��(V���?	r̴%�=�1�n�&6K�_��ˆ�=�6��Q� ��0�����%XĒ`0!W�b����[��G�Ə��=�5=&��
���pL��}��a/���!�b���H���/(�('�,d<��hϏ8�0�b�2�ڶ&dݧޛ�s@T�H+�$,t��2K��G�X�^EMcFv��d&2ۂ�eYM�8ZI7=In�D���7,�'\KXŐ��qa�6�^���V���.s�Z���t˜S}�����@��#�b ߖ���it?�ca�cp�_�D��"Q0�Ӏ�*�DE˴���qA g��@��a��Z��Jd`�d�X
����bP�W�4�����2�!H������c(��hS��+Z3q�U����� w@��n����\OY�LADٔ[��fQ �L�Q���OU�2->�ӅvvW����4�T�X�Ey�۵�F�  �Z�v��V^���Y{����Wsº�����
��xd~CP����_��o��%�y�J��E���s��t�Iv�'z͍���f7����,A,��/���Dd(�AA��Z߂~�<&�D�%5��<��|&a�����`��]۠�2޲�y�t~j<�9~��G�?��!�9�Aa����@(�L	�~���g��:7L�/�����u
<
R���
$x3���y��Vt22���KVy}j���-[��p�p�1�Ⱥ�{X��֮;2��<�kj�nU��=�=ϩ]�O�m`�f[�n�]#��Eg��������wXc*�����!������#E���	���z�B�&�C`-!gT<R1 ��5��>���;�$�9x�+^a�������L�=�8�ą�llv���\�M��#�o��j]�!2�r��R�����G�M��N�`3#��f��M���|��ށ怍MYo}�rJ(�E� �α��T3L8��K_�R�`�6�5���aY�z���\*[<o5ptʔ�n8,�V<�%���_�<��4��7�:�vf����>�-�3r� �+{��m��͙�O���3[�G�-�G��jj���P���d{hƼ�E�r�adF8�9�}���۷��-74y_���}�Z�t{_Z�u�Mo�2	��]`�Lf���X��h�Vv�5��cc��z��|�� Z���B�O1AM��!�������P��[�/n��-�#��=�	N�t��!�ʱXt�1���!!�b�ϳ��*��k-Oc�m@$��!$��eW �to���ޏv��ɺs��/��pZoI�4�lr|4}w�W����񬍏��/����DBXR��{3�\����,��莴Ӈ�w�Y}")��	� ���Ζ'��{��~�j�P'��C��/��,Yk|���kr���it$��);�3=�り��[�¿��7��u:N��{���`/������$O��g�����=��cNGcA���:�l��5���Kq��|��ڱ���Vڐ�)�zc��}��!��s
�}AG��-��`�}�L���y>b��#.�����0"�0B.������9��KC��]��{P��W�rn?�!��7�e�gX'S�j�6h͵����*�{+c�����~���dm*��]����G��~��Ie̜Y���=z\���G��O"�/��iC1�\��U�����{p�~Z�>zZ�s戮�?fc�۝�99Ѱ�;��W������^ ���[y�,S�L�{���66���$ͫ��t/ɣL
��(�t\#��N^��K�FQ��=���	.���l'	��K;(6����l�F�;�jW�ȚfRV�&�~����g0�>�\;㌳|--_���~�/�Z��[=�����z�pݢ���Kie������<+=��/�'�x��=i�֘�x��~���i�G���k��u{�K/�3�8�'��LJ0^%6q�#�8>�h��y��z �\&kQ��9F���0�s�(x/�|��f�tfs�����+�'E�8�<		љD�0d��#�,�ى���Dƙ���	2}�����"h.�c]����'�*g�9����SXO\O�qRP�!�JO��ݺ�lw$���k֬����:A�48ɡL�v�u_K�`�v��Q+�j�Z�CIy�%,�q�fV�U�
��u�s��DY!���R�>b~���M�/��j�aOm|����$�������Z��{vϝ��ӛ��W��5�`�,�+���6=����;�\�4�^�[�'ּ"�g�y��Y��v��e�n�d�c�����Aa��Z���i�sɲ۽{�v<7f�z�o��N;ͅ<�:mv�8)��đ�O�=c��G}����SP��^h��bzc��a(��"E6&�D�+:^��oi^��
�J(K��<���{��X4�!�ň��D4}�<���P�U����,&������,�邔�o��	�$^5���=��g���V�В�[�K�,K�g��O�ã�+	҉�,ڪ������d�����7����[*��wK�Sʼ�bm{�(��L#sK�Z#����#���_�`4�~ޒ����lI�'á���NL5l|l�x����/��b�y�a�=>əg���9`�����F=��Sltt��4��v;��c�ϱIP?bc��aU|a�	�vW���^���y�l�&y�{��]�轉r �o��o�k�q%��_~���D)�S�_����z�������S �K�ySB�	�L�
D^�ޏ�:#�^�}��)&��K�Y��)DhH�9����~
$G��5�ZP����5�,}��r����j(�e�A���-]���E�7�9� `hi��p�+4iY�4���\�w��6>9���@s�.���|{����o[���M�Y�E�N�sK'.�c�ȹ^}�7/c��/��7��G{ ]�|�z{����y1��Fmْ��s�6Wp?���SN����8RJ���;��x��"��^��zp	E��&�k����㫛6=n'��Q�  Iԝ?6e��
o��+��	�V� ��!������+^��g�@�cA��Dt��3ͭd��1��s��`},IA�����;���nd53g��&�R�c<� :�,���{#<����^S���XF� ��^��cnH���J�f�zbI���z����FV§�,ٵI�Z�ɾ2'Tp�����xF�M{?aɲ�~��oM�=̓�H��MP4��BL��t�������[�P\�Z����˿��EO)O��}��=��ԭ�uĞ���C���ڱǮ��kץgٲ�RSHG��/������?��O�|9�c�Gy��]s�=����L{K�]�¿Y��I��o��>�����b=�١���1�oƴq�&���O�p�|�^m^�
����GP\w�u�pp�	��A��c�wdg7�e���)��i�,Y�9FPJ����`+�+�N�U�Gʇ��U%�c^�6wL ����v�9��>�����=|c��{��v�c>�l���";e�J���,�Z���w��$�̂�N.�'y%����+��!��'��K���=�c�-s��R�J�����h�t\XK�����+�}��;�<��_�U���߁��xd�>�{�;����Xc�'Ň	�Ï�pX:��k}�<���#�<˕����ֻ��kiM4m��U��bMD�g�߳k�E/�{�RK��N�/��/fN�&βɫU��M��L<15Tw#�*���~�!*7��]�C?��ُ������U�)������o~�uW6�V|x	��M�yC�K(F�����G e�g�}U��0�!�!(F8�KxpN>ˉs����j� ��x&h15��"ry-}R|�+X�E]P��-���پ!�)}���\��,K�VYe`iV��<@\*W���=͖F��e{���k���L^t0��̋�5�I���l`pvڵM��Gg<%2�.��b�l��̅�#HX��G�I[X�R�j�����x.�:�H�7�CN�����d-M�-}O�^�ٞeH�B�]�¿ԍ��*����X�: ����g7�p'����崨�_ZN�C�)�Sw�Kբ��Ұ�y�L=�gV��63������{��`�j�� ��m���C�6�K6Y���ñ��?��O��uϐU-Z]�dp�^�7��ω�zXj��y�!�����*՟s�z,�qy��g	l��ܛ�N�.���k�\�"8�S2��jȒ�a�wZ}����R^A���t:o١���cɫ~����d�[�:hO<��Tyi�HR,��Z�]���\�YO$܋�U��F�9w{�x���퓶eێ,�ײd��h�;7Hs)��%�!N<�g�<���c����ەQ���	JY���+�{/�rqT�Ȓe��z��}�6[�r�mٱ����X��?MvO�<�Mأ�<��Q�O�Y}hZ��41#Vo���I�Q�vȊ[�{ܶl��欳�*�Rzy*�Y,,=6���h�(h�U��%�����C�YA�K/����R�S~A�?C�y��emɲV�%����0�����<G)��ȸ��T4N�:k
1���m�g!l����E0Od�Ha�}����׾6S@�v{S���ط��9$3U���-��cTbw����{�/�R��ozf��6����$,���t/O��q��$�К�q����K�+��4�7���j'�u*���i%H�^�mS3�k_��~����!��!�0(š����S	���^����d��x\�5�j������������gmbr�ο�,[vH2PmԞ���m����M�:)�4�?����W�>�,b��|�N8~��%����`��w�m~v�'bd1�J	����$�e�~�!�iXlR�{UeѼ���׼�5E/-"ea�qם�����w�/���b���nk�^�\�1cFA�Nn~dIȃY�A�J��>:���]*��f�!Ų!�.�Z�*8'�qxZS|E �q~��
���.���u��攋��4#�gF�TBV�ٰFS �j*F�ߔ���>�{d���`�Y�9��\��_~V�� u�/��H��V 1�+��d�`(�����v�/���7���������=H&�u�]^:f�-v���m�s������� O�֬]jûFl鲕����;�زQ{�)'y�J�����{�"ٞ�w�V�|`
���/�������ڹ��V�X�A��?�v�x��ȳ��5�竖���O{�����t����n!)���f�����G�f�����ۋE<:8vHX��M�9<2���Z�I��Z����I�߼�< ,��2�ʊ%H1��t}X���Y7���i���~,�s�<M���m
�CP�9�
�P6 K���R!���� �(2V�q��hgҔ؞`��d�QnA0L��GP6��J���������B��[@!R:3ɽr� �m\ż�H���Y��{��
 ���y��fB��Տ��Gp�q��e�t�HoH�߿�6=�ɦ&F��Y5�Om�dK�bkWeW\v^:~m�%{��-�u�D��c��V���0�)�΃�~�;��;���68�o�#%;��b��m�=�̟&�1�S;����/��ի�M07�ζ�~���{��%�\�A ��x�^np�7���H��3�����CPV0�1�X*���rW�f;�uZ���`I#�# �sqNA>���'��Pք���
^T^�M�`
�F�c|�-�׃����HB�\^zd�]�Cu��$�"b4��HT5U��,����e��T:�j�2ku�Y�	b��
���\��_��@��h͕ 17����+#����}
멼6�!�Q̳�#5d�w��;~�*k��ǜh��%v����Ș=��öb�!�b�Jמ�^t�u�zOv���w�{]R��ҵ``�|X��?���ߦ�\���j؏�3_�o|��m�в���^}�v�k^�Y�XC�w+gk�0, ������X�:��l@(�#��f0-66�~i�}pt�hl`6�\|��W�R�� ���H��Њx�b%|q.� C���C�V�`����Q�]���cbd��^QQ1B���׃�y{H1Q�2��}��z�R�S
��5������x��&-�
�ߖ��
�>]h7m�׳�Sn��f��?�{�
Q��r� �4�����9�������x�}~��󁒅�)
hdW)��*����y���=j+Vn������7$I']���G���F���/����v�=^�F��}�.~��*���MF�ʕ�=SʉA�����ܶ���.��O~I�*��<0�ԅ���pM�5��޻��	"�N�j2�l(�?�я��� Y���{.��U�����V7�F��o}�L��_�Ln�R0@��ɳֹ�{�O��;b���� ,tq��W�0G(`�5BT� %֮����`ۇ�r�b&�cP\��(^��W�ҹ�%%a�V?�60���<R�5@���D����Kmf0�C@y=�v\K���;�tx)�������f}�|�H�-r �=���Tn�09<(]�9�F~^$L);/�9^��o;���]l�Y�k�C������u#6�d��عծ��Z��G7gl�ь-V��3�X�¿�h:elddgf���&�s��o?��v{��G�\
�أ�v�N�e$�fvo��6{���{,�F�SD�����?�C��h������KH0x������_��p�YXjxp,�P�U��SO=5#t����'�E#�폘?CBRyZ��Ǆ)�}h�cP] �t>����G���,�I�F�JHIgA������>Q,JTV��;:��l�{�<���e ;���ؙ?�Y��Z���]�ᡒ��l��{��b|y�f?.|N�X�>�6bM$����I�p>���"���gV�����x��<w��7��	���o�=���u��?~��vc�ݲ�5��!�n����o۾��ȕ(��G���4�����7�X�¿U�N�ECg���W+W������2͎����h��@ڠ�b�U�z@ic0�X]*��q��;������)AE`"(������2 8�`a������M&�Q���+P+H�y��3��$P	�ך`�F0 x���q|��W0v�S+�22��Jb�7V������J̍TO�Ž3��4�P�PD=�{�k��_�F���t�l<��P*,��&� �C� g��A��R#h9{�����,���m�pD~�1��1xy��{���+	�������A����	ni�3��k_��?+�Eo՘nb��ݶcǮ�HH߅g�{x��T�̳Ƣ��GZ�Su���H��#ɵ���0=�:����i4������d�Q.��=���ܥF��D��44�����C��O��Ii0�0��#���M��N�'V��KL@��|�`�`�tB[X�k�軕���=�ǜ	A&*��?����x\k�vQ/���:��(�I�3ޟ(��B&+�*�C,��;dH �r�:����J9w
�%�Z>
�b����l���P�]�>?��`l���<���i6
%��(XS�\�6��9y/���l�|9+�9W2W��Ox6q9�}��H�s�4ʘ+Z"��K1���z`�(N
7�����=�����q��栘�A���G����"T��0XC��Qʆ�c+}e9S=�S��J��l�����d�Q|�+��E���z��ڸ����"b��lŅ"�7�\��K�D���E����BK�Pcq2Q�|sV�s:�>�wxE
^
�%h�������l��#��m(kz	d+�h���E�b09���e�k>�<�%)��ȥ㣱 ����ܷ�T�,�u�NA���	���me4�y_��tEPˍ�z1z���3V#.�>/�@7�̸�*<s*�:-�ޚv]{;b�yUڧĀ����@�����1��`��=�{�̣R����{��E/�{|go=���:Ӛ��6��?�y���aU��� �������>p�c[m4-�H-�9��mp�Z��d��ǾЖ�(��k�z�k#d�=�Ȣ�A���	�U�G-9x�U�E�by���Cשu��v�ɳ�x�X-�	%Pe���B��!ڦbU�������*��"�\D�z2��s9�`�}�&���aȋ�E�m�Iq�kjgHO�=���sYM����ڰg)�c�՜^uS�o��ٵ�bn�*Y���y���g3��s���]3g�*F�gV���_��{4g��sE�\Q��C@������r6�,G~�{�.J^l�.�@�p�v��mp>��N(`(��B`b�r���c"�Y�);ݫ��7�����b��u������0�O|�^�G���m.���:�_��`4����r�3zF������3|�*��8A8�Y�4AN�֕
�EA$�&!��w�N~9,�}ҋ�O<+hܫ��")
	J�U�b�n�2%1��IyZ���htXx����{�}�D͌*]��_aD�b��wQ?�)�U`����^������(�p�	�qi�,��YQ��ͭ@��T6%���*�Å`.�bC��Ҩ'X����õ��׮T�,��χ�/Z�P���8��hY*Q}%��g(�B0	�/���S���΋*M�0�CL��9kPP�2�uY������Py�����0�C�`�x�:��T`�)I{gEC��P�Vre�r$�cs)<�K���>JvblԿ��#��ƾ�[�x��5��PW�\�}�'�۾랻3je���3��"�.���yD�;����l��!o�y���G/�f�8��6�bD���m�շSC�J�Q�`�K	6Zp��TS�H6�m����h������X��}uǠ����Z����9����{#���|
�	�ݟ�{�C�A@$zqR"�^),	�s�~�o5fU�k@h��#HBВbGz�N��ۇ���w_	y1�$�4���nCumtm�l��~V�.�1R#���l�[]���%̹�Q���L+y�*q+�F2���^�c����X�¿���L?�g�5�.�Y��̔�� WPM�{��e9�/�_~Yb����f=��n�%��X�,/p�a�~-��u���L��r�|׎�UU�.s��9O�%Bϟ �,8��g�u�c�	�^��ye5*CT8�����$o	+��V6��:�X&b�ț��8ߍU�^��"�7]�O�S�A��P�N���X�VJ���,"�:���n�R�i/��k428�k5g�Y�	���3�� �C����V��a|1�C���ǿ�س��L	�1��o�/{�m[3=���L��5���Fĕf�`�j�ֺ,5Yڰlq�%P}��zo�XbX�.��r�^
v�M�0�F�L���k�cD�������� Ās'�R����}|��T�-*{�C�,oi#{GX3��n��_�ñ�,)�5)%� Vf0�ٯ��
Q��x��̫n�W�)�:8/�'�*,~h��>�=�r�6���a���O#�Ә��i�hOkϪ+\�w]�n�gX��sؓs�\ا��nf��T(ɐM�H�|�g`��|�X��h�S��j�K�F�/��P.qt�5�����V[xE����,#]�R� ��\ӔM��H@ĎO�4v��=]C'��=Yt�0�|C|�j�p����eD;��g��֊���1�1� n�Ź8V5���9��5[��,~,v?�FLYE ��T�?*w5v���X�3i���"���nR�P �:c�X������in����U��e�4��_�1�O�gQ.�Oĩ��L��֥�2
}]���u龳}���~n�Cy>�d���6�!��"_ �����@E�^���}(�P�fV�X����f�)�x�q'dV�Ĥ�G�mٚg�V����%�!+�����Z�F
c''��-vX�q�j�+`k�hQw~N���3a�^�NX�ҧ�PbP�G���GB!2g����PB�y��+K�90����a%_͵ܶ�έ��3W醨�Y#@�
��<�	U�Gx2��O��ד>��se�F>�=q�W\qEf�4��`�S������z) )�+�9w�~�扌d 73A��׭�ViZޅ�����K���~R�=8_�z���'��1���^�-҃Y'�p�y��g��@V�i��K�����
`��V�'C�4��7N5	��1�:'/y�K���3���)�:�&��d�y���'K^�	.&.��O>�j��~{��fcSD
!�[����`Y1�Ŭͤ���)dU����GL#Y��F���QK�G&	#*3)C	����!O#&��߅V 
�I�<"�F�Ne�
��^P"�G�\
E]��1>7�^BZ��V�̺&���:G������JT��!��2�״6���:�����9���z
ȫ%�Kq�n�[�Qݓ�Kk�כ-���u�s��j�+�"3$�5�2���G��^��N8�=ϥK�����n_?��Ńv������lyY�9�t>p3|���U�gVOQOG����|�7\��H�HL��f��V��&k��u�i��op��L:�~��~�7��_���\i\{���]Dlu&�Lc�4{�N7d�kX��%������Ɋ��YC����Z�Ŏ����N��ڬ�.��(����u-<�d������,AS���z��u%���6��/(2zCR���o��0^BK]���u�μ�V�iD���T�UDl����Dh'Z�b��we�f���lC��O����~ �uZ��W��(���!&���d`R���3�p�oȕv53��9�l����䦧�_�G7 �U"�P	t_Ǣ�y	�YI!�Ed�j|/��"��񤝫e\�qۼ#�j�e98X�ɴAN9�$[�f�O�����ª�P��K�����|�7ۿ��������^�Sة�	Pa�sI�P	C_MA�� ���1K! ^��C�G�j)���'�
�ٯ�r�3v��,x���_��(���Θ��/
�s�]�ys�L��zI ꘨e`Ȼ�=d#D�s�L*Qu�����y]�	����n/?�ZPRН���Q�1`�ƺ֩F����Y�KAc=��&
\x5Z����4��a��⾋Ɣ<���Ø@���կ����J¨lN��(�8͂$���ڵӖ,�����>�[�/|�Kɀ�ϖ-Yj��#��q_Ǣ������˽�����^��+��9�H���n���Y�W�\�=8O?�,��<X)Z+^�	D)<��#>���_����|�#^��f,���� ?�5��׆CyQ%/C�v(�'�9��~�(9~t/j΢���5����lV,,e��������Q�Œ��$ "�����qi.��z�h�Ȑ0��=�/Z�<�JR�1�'��R*�������R��bs�H�t��Z�E%�EZ�s��'[U+E�YJ^�+���q�6"�罠���@m�7%�̟����c�~�^ӱm<\0��z��ב��нy	���0������R���7�>	~��~��6nz�n�����;}n���=�<[��P'�,Y:h�~���_����^��A��v[�¿Ճ�59Q�`��]#v�1G����d}�U�?�arٶ�q��Yv
��/�ݞ|�q;�e�Y��RW_|�G5jg!bI���p!I����ۇ?�a{����3ZGmj�|�6��(l�}"@X�����k\�h�	o]�g��9Z�q=>��X�jT@�8�\	&Q��[B^TG0N~7z�Xx��6*�X/E����xu�*1���u�־p`�S�]T�A�-���y=Blj���C�3&�˜0W�a���=�X�ū 2ǣ�E!U��FC�q�Z�_/��@�+��(
���e�����'wq-Y���;�1��3'W"(��<m۶=�s�C�����h��=�y�k�A%��g��w���2I {n�3v˭?���m鐕�%{��_�5�����^w���V��UW������vNI��Ƣ����dc��\ȍ��N��m|�Qk�ǒ��O�t�UrL��o�޴�׶l��w��}�ݑ D�M(�#��F�W4<�dY�
|F7�׈L�N�!��M��T�b�Y���М�sa��@8F��x��
�,S�	�X$���*!#Ꟛ���D�I�="^�Z�RFX��	<:���l7�' K[ޒ���.��_�3w�F���������q��3��U0a���jq]��՝{���7�!�-4�5�>��Ϻ��� �8���q��<��Ig������ܙ�+�?�
�zQE�������o�o�q���\��1��?�>�[�y=��Rԭ�1{v�S�s�6[���zkmbr��Z��}�����ˮx��AA�u�v��?rJ�/�K�3&��Y�kIz��^nL$��u߽ގ>v��o8̞����L�?ɽ��)�oO�J��Э?�Ņ��ظ��8{j㦢 ����)�.���B�_����n�tz	8Q��^GFE�5�G�g)XJ��\��,>5���*����BB%$T�����e&�@4Eᘂn�#��`�ApR�k��vX��/4癝3ǡ����i�iw&�u+w���Y�\�փ:o���v*�^�J=(ʔ�����&R�������|�yWp;��el(�4>9QԧaD�c�F��@�ր��+Z���״�bn���]�J��v:xql�O!�F�<CFRr����oذ�~�#u���o*�;��Uo}�-Zb_��W=��o
k�b�z�+���+�mz�qk��؉돰'7>��~��F&_���-�����V;�S�_���Jo��hvx��@�������;��;�V�\�&��I_���u�G���6�`�)X�� [��1�,(K���kXO?���@*��𖷼�q>�,����?m?���E@/�ᴐz�N�Yt�8{W���B� ��,�����o˞��>�@R���^�Ғ��+!
S�uH�I���|�>�];-���k�gAO,�p�^Z�zL�L�Z�+��|�[���gd�Ǻ2���	B�������&6̹+�r�5��	2�ٹƤf*lV.5�&�������A��KVt	k_�����s�X�b)
����?���Z+���~��N㦮����<�����{ϝ��C�@J@�S@E�����T� ƭ�2h��� qd�	':DM< ��g6�A��+Ib��v�����R�d�?��S��-�m�&3�Y�T�R���L��h7�@X
Fbc��	�b�}�;�q� |�w�w��?�)��Ul ыJ7pd��������H�0J���	�$�)��<�J����ıD#J���P��I��@4��D.��1"�U�
���+���������;Q���>fbGVH�̙�ye�:� �ǅ�G9K�k��(
�v>g����g�W+X'*9-�W���fce־_���ݳ�{+�L�]O��:��ÿć~x��n��!��e�ā~YGxyt��|k�����m���y�!i�ҟ���N��O�s��=���o��VK�x]�\Ǣ��L_���0D��rˊ��Ov�����I�*-��!��X�C8��t�y�{�:��ƥ�'-ߨ�N]{�L��@Y�)��ׁ���
03x��4���V=�$P�(�)I	+}w��kr���B�\��b�;RW�rHiʒ�	Uz��+��>���6��ˡ5֔<��{���k� �
d���?� /�Y�����%����,�)gP� a�
���Q.�z9Nީ�J�=�L[6� �`���c��BI,��3�bє�u�O>n�F,@�%�� �D���-PE��O�S��4��i}Y����<:�ÿ������OL+s�)�ۈ����i�>����l��z�ȏ9f��t#�+K"�L���db}9������H�Q�H���l �"�;�3N����Z�!��|���ǚ�lv�HmhY�F��1�����Y��7R�$@�����R�n�SѱN��G^�8�ԘG!J�1����������6S�������P�q�ְU���yMA^�Q�C8��"��d2�R�z�/(���oֺ�ː�I�����?��X�)L)��-TF�c���$���O�q���-�׫^~�S�K��p��ۿ�A�w���M��w�y������>�o�!���[Cs��_s!�m՛S6���Z��rr �ג���2���Ĩ�5�!f��9�E/�ͺ�wgg3`~�a�j�a�;�OѶZ�VV����Ln��'m�ݾ!�p�$&M�*�t~YbJ�<� �"ZR���lC�����`���q 1��6	l,D-N����q�����=���c�^��V]A��y��"�^����%mJ1pH���+Ȅ��f������^�g.�_�M=7��
ݕ��uQ2���Aq��0ψ��=A2~e�j]�X��o8Ya{�F#�k����xĠ�����i�=͵�Ѿ�Rkv�L���mHc��{�s���W�ʧ���8X~�m���<;�XO��������X�3C�������,����lt��ɦ�|��>gcim�Tdh�
�&E2�\�¿٣����l���^y�����s^�lOۮ��l�����F�(��Z�R[����a[w�R��#I�[�8�2�#�KO,�E1(
�ن,���`U�W�_�;���}T���X���r��bPL�t�$KV�
���A��C�Kx�*����v�������n�M*�D�LP������υ�h��f=��1��
��2�A�1j )���`p>QL���QS�L�Ab�b���s����]��cnj��r�v�ry�z��0�-�=�N�n1�00�{���!}�!;�%��3���۞�F�φ��:��4�v�I�أ�lLϻ�pF_2F�3��w�O�&����;��9�i��g.8��$�WZ�@5�W#���:�t�?�g�Ɇsp)�v��.*0m&���l0�?��?م^XP�b���G{���ͯ`�\��%p�0�YE���>��f�9����H��s(���C�0F֢��V\��͓!�\�AyX/�>�5<��"��h���6?���$%X��P�e�� �,ƙ���A����H!w
"�Oтǻ�F��Z;����C���ľ�,��̚��o��33��o�s��&�^�9��3��潔@l���-oՍ��z�a)~�'��7���>��[�;e0�&Ӽ�\u��ܽ+}~�m����J�犲�f�d�Ye�^v�{�z�<{�F�����/�Z����'�BIf�;��~�n��&��5�Nx��:f�/͝���'7�3<n�rՎ8�(;��uv�y'���MǺb�p��^z�M7��"�gS1�K��B8W���Eb)0���lB9&����|�7C��K��{D����uQ�-o"R�Ua�XH1��x��l�wO O-��cEHE�L	��6��Y�M���3R��m	r��P�;��g�a�8����D&�����W1�"~��dp>�����`�2�*�9���i���b^�_s=)�Z����z^ܭ4͢oN���\���zT��*ʹ���
쿈�NRӿ�����\�h�����/
�ꫯ����ﴖ�<;��+��,	�I[��4۹}�y�i72��ɲ">s\20/����~�	�������n�G~�ȍ�t�N���*�¿�G�Y0Z��ot,���K�y�?�X{��׻u����/�ڵ�rNu�l�L�S����X�r�� ���o���_��c�4��;X߸���o��"�3\�cb�	A+,D0bY��,�IٿwW����/���<#a؂��6�%Z$�*�~�И����?
��Y�<�'��7T3ch�ƫ��x��3mB�<X���_u��.R�,e�
�g�x�j��8֥�-1+���3��^�?�x�.�����Ox�bŚFsabE���B��B�%��J���L�dk[sR}�ݾG�K��BŖF+�q�Y){���m���Sݽ�^^����~eE�&`�}�_�ߏS�eyƬk%H*7C�c�Ĺ�/�ܾ��>�ev�y/�����)o��x����������lȊ�ױ�/�>�wı��Ѧ��g>�Y����� �v�����8*���6:Fᬺm߾���o�օ��ZL�����x���������.� ѧ>�)_���]��ψPL��Ŧ������ fHH��8� A�(PX��s��糲U�AHΏb�R���
���:�%���M���D�,T�AX�|��2�D%�
�1)�z��_��_�k/%ſ*PƘ�k-v��Ǫu�kS��
�	$�.a�3D)�9X�Ϫ�C�T�����JaP���_��`!�i��>A�F�!���"��`��H��9�%T�NtL�@5��`�:�t�&.������d��Y�ֱ��ã��̳ٺ�r���2�;STޑ�zŹx�=O����\��x�rX �7q�o��^%��K.��Q�s�)g�`�LN��̵>�����{F��j�k��V��_Gg@�QY����W�CP_p�Ey�⩂~���?�1woQ�E4K9Y0X����Q�෾�-�.��B/�@�@��
D�E��3,y0,BY�
؉��*E	E�D�Q�/����|��F��.=��r�=�C�"����@
�r��'b�,4��7j̑� L@����ΪT�EtI��Z�ipN�s�)���2�J��9�[��*!+[qU�d�c+P��c��cL`�!E�ʶܻ����c���x/�"&҈�(�]p~��'ltx�=���6�kGz�n�[��R�"@#W�<�,�Q돷#�8�cqO'��^zzs�-͗,�93�=�,�'��X����Po��@�-�l1��s�v�w��x��_�m���a�g񙆓���k�X��sN��?�Yͥ��q��/u���d��M�\饎�e�Ъm|j�mݶݾ���x���k4�%0>�Sݙ�����
�J(�E#�x��21�*( b��JP0*-�6�'˓E�LD%)H(]TQ����'�������#��Y"A�� )$��n���V(�eM�_�X�!���w�k�Ϝ��{|���3a�#`e�G�q���C�Q"�N����wz%��x��ށ��4Шp����5�Dzyg�\u}�A�ɱQ+7�WI�F_��+�Y�MU�-�D���X�]J
#c�4�mE��h�s)�/+�s~��l��r�AG�^�L���y��
2�JwH���o�F�G���xR����p���y*s��N�j#���x����e��RT�^�+YU$`d�{˃+�mg�wʭd�!�x��;�g�UC�e�C�^u�U�(O;�4�H���T���&�5r���| )��X�vK�ɢs#���d��'���|*=��Q�?�ѹ7�AX��? �]V��V�zY��k�J�Z�~��`���)� L^������)oa��TyS��UDN�[q<[�?XW*/�h�9��b�sC(���'��@&�kdl���wHA�
*l���E���~4�C�.���%i�٤��[�}W�fΓ���̠R��M���ʜ���{ �v����6��=���J@g>�|�W�*&�{docpѷ� �bzzf�ڱ?y��2�3Y�6=�%�S�!����݋�S{h�sT���g.̸R�t`Z��m�ˈuWD�t�%�_�k�� ���`���`�F<�k`�I������E���'?�Iߔ�A�p��?~-W,�����W�v&�)���,PY���c��|4�N� ת�c���`�^\R�����p�E�YpLE�8�0Q#m�K s�Yo�f��|.�iމw���L#�de%�u��iK��ol�+v�0�N\~=o�yQ�D�7oRק����T�X��x����p�u�0o��$�T�GU,X�s�%�e��X7F��l ��{s[�)7�j�	�d�I�yyh��@溪bB�AmdD�����y}��_�}N�7���������̟�nȐf��J_�&��V�Oϴ�ɣ��~�ûlp(y����ʔ 6��F�$���&K���6Z�"�~�E���f��d��m�z���K�1���R&,����� e! (���O���-n�IH�d��h�h}Ja��#��%oɲT0W�Q�'z�+�:f�"�x�AB���E� �K����0R�N�
��F0�@�R�Q)1
Aל�ZKi)�b&���<������H�a0�7��%�5=	 ֔�y�����l#�1⻕�a�r���I!���g#�-r���X\�ۂ�Ӝ�f�Y�i�%%�%~a�;%t2p}U��t~�Ԫ��!*�8�W^��ɑ<!ŋX׼Ϗg�潒�HX@`��dՍ��'m`{��J�V�Z���I(Zg2L���Қ�� ��}5�x���du��Cm�ܵ,{i��H��Rő4��0�O����[9_p�^��w�>������M�{d�S�c�,�����˳keMŠ��T HG�B��x��rs�Yd[%�D�dh�r܇(�x*׀`'\�d�q�QF��D��7�hΫz4�.bYDG*cy��[FgPS��C}�f�u3�ۿ��΍����s����<+�*q� ����ׯ/�S�]�j��bs
&� �G��<)��R"XΚq6K~OJ��[�E\ks�,b,"Χ��2�ߨ߇ ���N�C�VL��<MQm�3�۩�1���<��|��6F��~��Y�H}���+�$x�PQ��<��QfK���0�־A��\��G^�d��3{�g���y������_,�i*��^|��2�a����^_0L',"�}ڵ�r������z,��c�,LYw�?`���>���x�*� �BP����[��#�&��,J���Hu�`�}�m�y�G�x�l��1"J�P̭�%�n���@���8V����͛zK��,TxO��I�L��Qָ�4t����Cl.�A�~���$�8�g*�=�f#)����ߏP�{E�¸)&#o&��ϕ���܇��R�ϲ���D�p~]��}���o~ӫ���?�q��C?���eĐ��׬C�劯!�F�}��1z����ح�0�j@��EL9��큪�k���/��/�ܲC��h���;d9��Դ���zt�&�F<9v������mL�(j�oh��Q�H���΋�#.f�
��&P�Y׫�$�#g_�X�F�'���{���s&�G���*X-���P�^��+Y[H��!K�&^��Y�xK(�X�ZZ��-?x(O�q*)A^S�G,I0SPV����-Ԑ��<f�S4�͖�"���ͽ���*�`����-'k�Y�y��5���%zp{��kDa��%(��vT�Z�>�`1����6<�*��Zӕ���j�i,k��f2�H���HY��}/�r`F��e){������Y<\�@PDw�!�u^4%ܦg��R�����9GW<ZȲ��Q��b���$���~���K(�]�ML:k��_���;��$�:�[c�}_�sӼ�p��7�SA���@y�E���yw>/A"��WF�^cJTQi���s�j:�֞����4�߹���ӳ�wLcy%�G�n=�z#=���*"��6K�P�-*W�,�w�`�����<:��)���Bs~���x��PL��D�P��zS��s�[ƙ���dzɍ�"�n�1�:iN��|��¿���5���6y�	(հ�ZY<�'�]�/��z����fV�g�D	�J�m1���[�i"�:V,�SP�S��'���}ˊτW5�κ?1o�㗒yH�JTN��,��Y�m����ڟ�=�OV���b���)�d1���O|��1�S<��D�%�y���He��;��G'$ة����^�������b�u�T��'w`b�&Y��$k�{�f]�X_{&y1��z#�1�ǲ� � ��ڂ�<�k��;h>y�R��baC`��@�xn������9�Cc/0�����F/2����,��=���X�¿�m�6��$,�k?:U��m¶թ��6Fw�7c\0b�t
�ο�ń�4�C����F^�������5�f�ĲuQ�IE���_�F+��F�ә{=�,�Ҷ�ע��:b#��<���&�'���a�#�FU�-�!VL�W��(/NTP�(����� ����wu
���9у/L� d��Ne;�!ť� \1��S6����,߱d=[s2��	�	/�W�Z�!�\[�j�-]�̃��t<����.�O��ؒ�����Plѧ�*%�h�id�Ǖ8D��g0t��)���d�������`�9`���E�pl������/{���DV�m鲥>�Ln?cc�6�d���Es���
�B6�Ц-0�N�W>.Ta�L	�t���(�'�vۣIVP�s�⎐N���Y�A�N��Xݓ����+u!GTz��Fe�n��4���M"B�����.��~XX�w8�o�D��9����w���{^ÇzD�b�������\���y]kGA�R��	r�	�ס:R
x�� 
 S���p����jVճ����o��=�P�m�>b�G��i�
��*�G������|Kqʛ�BVv;����$����iLi������u�o$'��%�<1��o��\����y��'-+����ױ�k�n���vZ��	(}�}�km��徙֮]�Ʀ���f��[�~��<-	�G6&�@�տqkK�D���f�p����v�
���`m���i���xq(����"�9"]0ޓ���y�qn�:���v��y�}����O�J�"�M�﨣��F��w�^��~�Cr��,?������sX��\s��7��M��W����_��_�b@���}��zPԮ!�Tɂ�����*�G������5RD��5�C�9+�	��O@�G]޴v��p��,�JF��9y�q���=mKl�r[Z���J��)����$���MO�j=�G=��b?�'Avj�Ɉ,��
�F�q�Y���>���m��?X��%Mf�_�'�hc��?Psh��j7��ױ�?��f7�VGI���s��n^��Wم���d�(�sءk�g��)�'�z�]w�u�%�41��o����o61�෽�mnݱX���/yIg5[S@uY�>_��~�~7!*7�xV��18�4|-v�K���������{ /�	9�����VR�o,�D�����:2	d����C� k-��ɉiMTp�D�Ku�ԴE��=^\$ŦGy�8< 	Ш���5����E����iT��?���(�����n�����.U2�%�Ջ��:5s��U���k�:L�\y�u���-�\��ǾZ��w�@~����,bE|�w��C=���_b�]�^�EJ�ܛo�E��=���v]�����l��n[~��=�ȝ�>�~ g�v��=`䙝Y��$�)u�[�f�x�Ŷ|�R�ԎO��&=�ӯ[Ln��I8�����#�����޸%R����]�S���?���`_��ל��~�Wx!1<	Tc1<R+ƓO>�/�>�����3���ҏ
����	��Q����+�O�����;����R��I ���תe���Tc6���j,��CQ����Vj/����}vֲ���l���:)q<��K(&��}}.*o)J�n���uia=�n��s��݉-��-�J:n~l�^_�)k�WD��9�6�VS���8i����������#��j����'�3��ח��d8��H���E��e�'�,Kط<�E/�K=`�r��V�q71:n�sn�'}�L=�ܳ������m��<kU:yy��zꙶ����C׮�+��F�=��;��IF���>�9��N��3N;���^{��Ǽ\0�T�+����\d*�L��)���,J��~�}��fk6�Q)���
�"I��Ijg�3Z��<�x�#6.n~6�m4Y�p�I�X,�o|cZ���
.��`��Nq�9)g%�}�"svr<���z�Q�����VI����}���I�ޣ3���l\��{t,�4~?�WJ�)�K�)��g�3������͘k�ǈ��ێ��Ȭs�w��y�������q��z������V��hbZ�d�o�fO<�m۲�1�ի��I'��%����)��d���a���g��c�G@{��V���\�d�Vl��ەW��IcjĞM����~b?�$ؓ�54�'|��m����9�BW e,e5ؖŀ�Ǌ�aA�z�E ��&j��I��5im�[^�="_XV�g�Q��6�P;:�Pu2p4�	ୈ�a��4��HG���y�+/A�wI��r(Ы2\ץ��=<)���p_L��1�O�ڪ���;h�e��[bj����b��mt���^�!Gk�!��������M�~��ݓ���^
ts�>^�k^�;��#lb|��Fw�/��~�������l	r&I����y�A;����QGW���w������.��|��>ϑκ�c�+u����Sq���g����u62�ê��my��$䟱�]f}G��� ��:"�w�����9�W��J������g�E��br�>��F����{�x���}���*���;�Y����k�+�$'a��6T�+6c���덂Q���*9��-��_��L�+����P�G���"��9aD�"���1^2�2���|�
�1��n���(���X]���2�w�����GM}�za�0x�r���w��&���3s���gG)q�?�"Y�q._����*▍���g�d)_�k�8��f N�y�+_�kO_y����?�coV�o�Ϳ�?��?񹈙����?:6l����Ϟ��H��#���Y�i�9�A�뮿�N=�,;�����Î�N8�6w��	!���;ow�!����j'�t����X5�?��F[�jȎ?�����4�c��J�W�1۾c��%�Ɗ�k�a"�ُ% ������C�1���C#0\�ˢo�34]��t�c�AZm']��Ϊ����<*���������Z�^fA�H����6��"]K�������X�y	��>/ap����e0ڨ�
}�=�s�;���E��k@��;�����;�)ԧ e��4's����#C�f�3	o�S�����\�����^c��#���:�,�����!u�t�MN � 6��u~�9�V�f?l�=ro�)[�n��?��F�G}O��Q����ϭ6<2a?���X�'�֭q"
��=�Yi�y�^��X��d��v�y��iR[^5���n�7��r[��{k���"ob�N�ɢ�8E�Jε���<xKa-�9����*ңW�EQ,7���p8a�ެ��Xp���ٽ�����}s�M0:��3����R@ΌH���Y݆�U��N�������)�/�P���ΊMlP�*��y��*�8��ň���ǡ��ӈ5�E��#�TВ�'�C��b{	�={�uf
 �N9[ڿ�S$�u�?�;�:����)��X�|'xM`�[�pσܗd�2[�z�M���FQ�u/�����a�Q�u�s���`��w�{lx���v���E�����w!\��g�ޘ��ݝ}�����NZ���`j4�=Ѣ\��-O=h#o��/��{׻��X�� Y X}�����z�j�k�GKMp��ǋ�'��%�c�_���V6�h�6#ŲS�+�+�!�XL���*�|����U�}a����0��RL���k�+Ll�Q�C
4�q%�s!.
���	�+r�9��I	h�u����B�뭲[�e{aÜ�q��}W_}�{��f���|�����ݣړ!�9�{��s�l������MM&�0>�{a��¬zg9���z��f��
�x¿xT{�����{��ղK�V��*�_�����¤���P�ȳ--���
�����eu���{�m_�e��K� "mADE�b�h���-&Q�����"��b�-�`��BD�FT�" ҋtv�������|��~�9��{������ܳ\�ַ>�yN���]�AY�x��%/	��������,���k��qՒQ�>N-��U.���f��Y�x-C�(N��9>�#_%��lk���bm�m��R�f}e=�l��g]D�)t��8�����|�]���g��X���/�:�|�Qh))JUH���<ήJz�ĸ�X��u v�׫�<某��c`YW��؅�[#��i�9~:xp�VdG�.}� �>�>ѧh>*l�e�;4`sk��q8�}����Ͻ�֮���2d���� ���zu)^���oV�':0X�n�`X�|��$�H1�É- �r����� �F-6��A�bn�\~�_X��$6�`}��Q֐�?Gǘ�^i�öYub[�2�═��Aơ8h 9.�Hʿ��|�X� (�FP�V��H|��{�j"��~А~���x���V����7|ܾ�8tͲB.tL�`g<LQ5�L��;5�,���h#[�<�s��ʿ���a��Yk�=eH���\�(��?�nr�c�Q�hw��.ŕyvg�5�7l�Du�n$���Y�/�"�����X��<�Jޑ�nl���۲�J�2�eO��)���wo���w�)ny6]�W�8�)���1�0��+R�ʩ�|�{ʽ)�#���I��O���]�7{�����E�Ѣ^5R7�L2X��e�s��$�|�IV���Qԋ�o�L{�4��e�����ްt�n�)8���kV?֬Ò�W�9�^����%�Cm�3<��6������������@ ^�e�h�Ǡ���/FȂV�2mi�T�b�J���bT�H@_!�H�Gh��RӾ&J|XM�Q�y�b�",�u���.�-PW�����`R����V=�Hx�I���Q9/���JX�t����[n�3t��y�Q�T��r�%��:�[�떱��X�^�[���7|���8&�tW�.�v�����~�oX*ЬZ��/n����Ï�vTN����7��Ƴ8w�q9}��3Xy�ќ�MqKK�e	ζ�egY��|$P���լ<��I��S��OsǗ�����>'*��������|�0��.�̌=��>��]tQd�6�o��݌qu���¦�=Hݑ��m Ϙ����;<�ȣ����]����"�2�z�O�4 |7��J�և��7G��~�3�mrg��w���M�{�N��`�5{n8ꨧ���=.,^�gN?@?OY���s����Y��E�j����7�y��=�4)ShK[���p����(#�Q�=��l�Դ--,�5����WD�8�a����m�<(�����%��P;$��u�3CT/a�=��fox������j�8��#�	+��:�ظ�u����?����R��"��dfZ��&an
��/*�+���85�}��ap�?�ߡa���	kW�
�7�7��yX򥳣'�^Eϓ*K�����0��2@��Q�*���}p{P�L�|M��a��2��4�k�TO��C�7����a�\���e3�o�6jz��Z���`�	ƭ�>V?�"���+W�Pm>�⇹_���I"�s�!����懧���s@��Ca�ڧ,��v�,�=�[�(���Y�B�7�䧡�ws�M�Im�����vا(��	�	��VC�˾���j�S��SN��˼��¬��aϐ��VK�x��|�;V��V���e��x��h�nv�@�ɏ~�c��a��Z�CP(�n��۲������M-��q}�-ʈ�K�N{�*�s�����{J��n��p�Yg����}�d��#�/E_@��
B'�+�/�z
�^t�������9+,�u�%�}�'�,�������_�첼��r$�-���E^�&���/̒QI5m���L����ζm蝑Z-�6eE_�r�e�a�k�+,_��W��>��O�M��T+�_��B��@��mT+����g>q�rN����ծ[���%�r���4�<��wɋhDR+	kO�,KO	6_il�`����%?��U�V@�?0ʒ�_.�x�ڟ���U��:0����y�v���(9��Q��Ch����E����?/��� ~��*DЧ0�{(���;�x���g��Hݠ}P��_�����|.�J�'�]ͳnf �:�R9>~�!�ED�o�`�P��}����eM��R��c}�N��4���~�㟲���^�|O��Ю���#��!%)k��MB��e,K��O�h\�"b��7�#̂��0�ꈕ�+6=d+
�}��TV�k�b-�����yN�f��G��U����
A���3���n+�&������O����?G_d�Ϫ�):��/���i2E�U��v�IR����i���f� �{O-"cf"�r�?�A]�=B�_��W�k����eFY�E�<?��,3\{�V�s��#?��T����f,�_�Ѷ����0��=���n��PTG���R��&��o��P7�6����yG��޻�W��+��s��i�Q��C�AT�°H	8 7S��$�E� ��J���ۙ%�dmx�6��-B@=�M~OG��X4"
�RĈ&����j�,OO�e�����h'���.ޞ"[���5LjI�GA����������&MGƃ����i���2N��E�k3kV�Q�Jɐ+i�r�r����W��($�y��mA96%w5�՜E0l��/�B�&�\��%�7���1�ph��~sK�H�:���>k�H>Č��j3�ᶞ��?U��9�����P����z:�j)q[�,�tp*$ �k�z�ue�{��&Fb�t��(�d7���<�y ��+�q�WGY�ry}�F��� =7�?��s��t��X��u�v�U#j
�� F�LDj���m�r����H,
o(t�SnO���UDcK�Y�'B҈:z2E���;�1����KII���@eT�o�q$�~�9�OCh5Q�0�<�@��H��QJ�s�/H�[� ���/�c�h/U�(s����z���������>���)���
���>M8;\Q�&WR�,��lT϶�,�� �b���k!�|�;��c-fċ��ѷ����',E��1���[�Z�|!J���X�s.B�t=4h�Y�:&Ÿ5���h��=T�������Gu�X�;���Sr���)���=S�xD�!�U�Y�IcE`_M>٢1�á$;���б+��ΈC��ԒQ�D��'��W�u�Um��)<�n~1��8 y�˅�Ȱ5��f�%BX%#�K�~���=X�J
�n��M��Dj��V�K�����?KWm�MT6��ь��U]����\��)�	�w�+m͗)�Q4ΙE^�p˾� �$at�W�}*iE�h{���qkI=e"��m&
/�2%�\��EMqT�Y+�;�[�PQ�Mݴ��L�z(sQR+�9ޘ��-诮k�/�m1f+�w���dS6{oᘸ�,TB� >�篙Oו,�&o��y�	�Q(��s��)�Сs�O�_����2gNOn�#D4��Bm7k#y4XN�Q�/��C�1�a�V�6h��e_�J=�7��Zr1�0)%P+��>?���)�jV�7W7��7V�Z�u����4T���|����{�M��=��1��n6�=)"OC�WT�Ÿ���0��l-�E*/�,�re�v�0٬ �os��$����>,�d<��Aw����U�E/�!�@��C��X ���/}I�m��ro��]}��Vs���dJ=��Ʈ���/�xw�dd�"R� �'bl���$2BX��x��DSH/��-�7.�o{z�,�P�s�m�W�(�]�R��!:�d�y%M�p�J�J0d��\�aK�A�����~�s��y=���<�տ�Y����@۰c��3���Ot	B<Ǹ$�c��p��Q����b�����n��-��1�T4��șlM�k�B8�evi�x|�+��T��RMR�w���B�#d��q�$�uHť�b}�"�h���Ȫ'�@� cJ�ʾA���d��>~��*̼�9����5�8���d+���IG�*�5�&���Ƣ΅��k1�$�ܟGQ|��������x�5؂8,�Kc0����馪[ �a�m
LʉU�1G;;���\(��P�\�|LZ���u�!�ƿ���Q)���l
AC��\JW쁡T)��;�)r�W.���(&��A��H�=�C���{p4����h������g<>��̍�&��8Z� P��j��eU�I�s
x9��;��H���9)t)r>�&�硲*���#
=�O���X�"ߏ���T�E&[��ĸ�CD��*��h�Z��
z��-T�̪/%#�Gڽ� 3J5����ǩ=V	��~��&��[����\�W�Q�y������5)Z��������aJ�T����E8��Uμkiv���~���7�@�����J��9�ƴ;�o+2��x�::+Yf�ìl� pߌ�;k� 7Tqq���F��7B?�Z#񿑞�ږb�����|%<^��5�h �M*���B�c�R��������H��EM��\�{�"�7����;�;O���;�֌R:;���x�o��!����iҎ����g�C���Pv�Vݛ��g���c��E�wnM�y0�chA�}�g&�����3W�N���ם����`�ީea+Bf�yXI5A}}t��2�s<a�i�����z�IM�3���L)[��m�H�T�)e0�5��"@
E�SL�m�_�BXF%�)�k�c��L��SD~x��d'���O�z�a���m"��V�7c�X�_罴����}K��z'��|��exoK�TA��[�mlb�ް��'=J�x�޷���ֽ�tY�=5��\�3�֊�(?'u���|�ӣ������ȡ�S��Q��T�F������Z�q�CU�$��y�Y3iy�!����o��Ψ����)nx޼���a�:KΤ��(aҹ����M��h�7JVB,������ ��/Z�>f_T�� ��%哽�8�9mmry[$O��J9W�G��U�x��=�x��<9-�x
1�Z��S�L�xX�{=�Z��S��)q�v��&)�V�I����"Aj�a���[�$)%�v��a���c�h1U�I�� 2\��&��h�VO�q�Q����PV璵��r��y����s-,M(��`s�V����:`�A�����,�ߕ�����p�QG��sS8]�\J�}~}˯��<��Us"J@M�y��3��{��lq Aʊ��_n0Pߔ��58<���@�b_֢�W96S`�|����~���� te�q}szYt�WŅu��3���
!�d���������d���־��V�1�R��� �c?��f�7���crkI��b���?����j�	��� �[��ih�/������B�Y/*����ہh��K)�)��;��}�1F�ĢE�æMBGg�l�y����52+J�X�K��a��/^b<�rw�m�d�v�a�����y�T�9�~��������o;��W�J��q���w���ۢ�"��|ޚ�R����)Z��f��Dy���yL�"�u�$W�����.Y��&�S<~"��H�z�/U���@D?,�e����{P��M��D����8/�4�y`��+�YN�o-��A��-��Uua7�l���x}QS�1T�e���3�����~�Zu+�
�y���c�1Ѐ�)��y�q����~��[r��$U/'�iXq�I3��Be�%K��A� ���AR��eɀ%{W�^c݆@[tvw�=�\�X�$�_0�������������{��^'�/pMn��_�j���Q"�R���/���(���b���=yWq���B�ޢ-�#��믿>�
����B0���U���+o#���xg��Gl�	��ҡb\�;�L��E��Uա��>g�y�s��1�W���>�_g�>���=��¶���q��?�����=蛡t J�����'>�<Q�y�E(���;#r���[��H�QI�D�澰ے]ü�¢Ż�����ʹw���R��k��^������J�ț^��4gx�s�-�y�TNK�~�âӢ��O{z�k�ea���V���f��C�A��.}<�ce��DV���6@��XZE_T~>\����mg�Z����?�c�¾Ta-*
�;-@=	r�P���*>?��#I4&fb��6�B�\���?F=lUU�f[%��,a τ���%����w-(|?��s�T�2?-����u��`h�m?~_%�Ѝ�������*��g?ks�¿׾���P�P?|򓟴�#T�ƴy<���#?�@'��=em��֭��"�i���Jٶɼ��l�΄�ǳ�O{��L�ɝ�g\�l�p�����&�|�/¯o��ݐY�������=�����p��Ǆ�p��X �|�t�bWEA�k���lٲ|" �JV�౎���'��mU�H�6����,l!���F��b�ɡ��呕�a��}�"=��������~-�o��|��0ط9��prȰ��Hj!-yL!��rHߏvr�c���g�����և/~����LY11��ΒmC���ů;���SO��:8���^���/��b[���7m;�9A�������@�>��G�7�����'���=��~����"�(�:!�C����|{z�V�a3^�w���`�شV���n��e(*�êU����-���a��e��]�f]�ߟ�8�\�.�}�����'[G/�w`аYYY����c� c(yؖ�+R��OwԶ�jR�*#�oB��;�p��z*�4�)������p%+�V�U#�z)q��0̖����]��C��ې0�1E8������'yY\~�������ֳ#�0.ޠ8���z�E
LCu0��ۻ�=��*�a�����Ɯ���S�ׇ˿�p�	��7d�'�n���p�]wY$b[��i���&E^p�E݃��|�����/¼��a߽w���#a��}��b��֮[���p�?	���ߔ; �fbrr� u#�+ĀO�]A�����}�(i+�)-�e���"�C�������~7S�s�N�<GOs`CV��5� �~��hd%��Y��?I�Y�U[J�Bt�kr/��HG;�C�����cm���߹"�wιa����&Z�ᔓ�̛֬~*=�x�4*UxҊ������Q�$�a��Y��:�?@+�p��>�W?�fU�я�.�=��2�p���L{�J�#~��K��i�{`s_�;�ۚ*<�όx~ظ�'fq�rW6[l���u�6G��Gm�?�\A|��Y�SLX�
��'b5!�|�H[��-�l��hY�SY��y� ��X�a�0�ը���8��Ba%��b)U�fϙ�'�ߓ~/.���^EV�x�V@�/�
�^w�u����N���뫮���,���^>���Q � @��#�S.U��o�i�c�°�^KB��ު1 ���\w��`X�p~����-w�{����@B�ΪUOm�M{�_
�M��;��sٞH�C�#��0��qY�������\�a[X�<'	,�/��~�����;��=��!1��f1`��җ�d��3�I�D�ôe��p�J��h��^1׎DB5�bHJJ9�laӭtf�
��BZJ-yC1Z�n� �؜ΰ��Ѝ�T��I� ã�?���B<��Wq!�hFZ���O��-���7�l�n�Wy�w2�V�ZV=�xX�����t��l������T�2n�Zm�E@����L/�0����c�3Ꙕ��p�7K����ņu�CgY��MiqqʤV�6��$q�2B����� |F#x��|�.����t5e����
�Lm�W}�#CuYM�=�C<��"�r�`dl4./�åa�XH͈ޔ�5\F\ �� �M
?QØ�@�P�ƅa|��;�y^�2��z����s�����/��'�c��) Taz�CwO�u�d΍%�nI�4�
�Sփv�k�L���o&)?�4������Z���S���:-�M���v�OWGw�<0��ss�ӀQӖ����4/ݼ�+�s�9���~`�_����芧��֖����K�no�<�4�b����Q��r<�h�1��D�G?6[�5*�ٶ��u;O2�>)e��Z�	`��::��M�_砤����@;���Ë��E���/�x��q$��k���4�+c �Q��e �}�O<�.�E�ڊ�Aӿ�=��Pn�R����`G+{����ʺ6̟7� Vs,�?��tǬ8@;�������M�;��I� �"�Í�"O��$�2 (���#�?���?��?�/|����W��/(���-����S��{�.���6<)Z�C����V��k�eo��������'�������2ۢ�j��;j/(+%��E��*tQ�y���z.�����WCw>#�G���X?ߡ0�a�
ݺ��tu϶�J�fx�����5{j����ua�^;�6�gI���%�R���C女p���+��nV)u�q�psX�vSXs�TI����6�n��=b7�?�b�<n��ִR����t���Ȩ�;�n�.��_�o�}�C��N+\$���e�cnˎ�ɄZ'�TQ���(i��0	�t'�P����ڐ%q��*Y��?�i��xF���O	��`t!�d@���.� Ý$Y�_=Ҝ��-�fT�:�֦�����a}X�~]� \�g����x��C��Y��N4 ���MF�F����	�6�
�V�����{-�#���;�7���W�5�����Īա��k���ƀ�����B[�]K�i��s��VD���p�aO��zsX�a��*����[騄����~����ͻ��s�N$ox�����jx �@l����g�"�EEBB���Ԗ����5/یs�_u���������uM��RW��U�P5mi���j�����\��_���Z�v���-�V�%�<1�j�ق�!v�����I�U��9�<]�O�����{�Wx�oSX�iM6�g���U�[I�ݬ�粽�I���Z>�߰1�u�=F):���d�S�eȚ>몃�?�C³�����Ǎ��'J����3kd8����Z��QO;&�Ǟ����k�F����mA�g=�n����j� H�PZ~���t����-h�Xpmi˶�o���� ��w������y}���z���ʯ���Q;{�_�|��&(o�=*��>�ݴ�8��_g��W(��ܠR��\H��/|���^�2��R�c]�$1��0�|�~��������t���/<����xU2~��v[N{�s��
s�.�c�����]w�6�t��;c��5���T��!�w�WZL~Y\�I�{���|�>�Ʀ��G2g��ea>���ub ��e�p�~���VOa��
�ָ}(�W���:5ߞ�(�����J_O�M7�d�1ա����(��� ���O�H� Ҿ���U��J�����i��R�导� ��9�=�г�q�f�!`���A�0���9>u���W_}u�m�Ea�ys��y���f͞V�z2��m�r���|�5����7��^{ì�9���U���o&iB'����������a�����a��9T�����oF��~�j��FTra@��+v��;��U�<h-�do[vv���
w�[U���o����r����zܨ��0~r�?U��ߛ]�z3�f����z�*�J[7��,���
�b���׿��]�O����(~y@ZL��^~��-�=k^\ ������@�ي�2cq���QGt�u��{��U+-<T�3��m���q���Zޘ�%��/~�?����7�����q��W��6���ׄ��+�巈���������fx���;�>������28���w;�Iy[ڲ�ģ{<���jCi�ݼӮ����m�$���y��6��gaTY\
`Ͱ��l;�W!��"�c~����I'�d�Y��	�b�Q�N��������O<eq'|�;��:t�;(b�i����On��y����S��*�^�7+�R���m��fϝg�W^n�����u���LY6i��?��n�:(-'��!]$�����>����f�q �/\`!{�ψ~�c3,0a _�5=`۲}e���L(��̘������@�u�E��8\�`��vBj�S�UΊW;�ݲc2�Y��r�c�D2t-~��`��>I���_���l���MA'9�o|�F��^Q徘z�B����|�*�n8萃��˖[�?�G'<��#�E`4��\�6ܗ�3�B 0s;y5asey�jg�ǒ������X7��?�x6,2���B�=����W�j�\F�O����
�����G\�mi��*��0��ϕ���	[�V����%�����{.F���O�f��Y�[��A�VT��OA�5x.�³4jBA���O�~�к�{�F� �
���Y���Z����O�G{4k��:+{h�����z���xB�X��}��]�5�`-tf�a�q�ש�Q�d
��J�!i�!�Ց���^X��/�� $9������e��V��(`[L�V�}�X�FZ��w~K�@�������	g!�<��/�	���5�暩�����:�*�B*���{�"X`% ���~};P��HH�}�mn{J����3�Z�V���Xv���ζR��Ŏ�ي%tS��
QV�(�T�b�'�ݡLq��ϊ���H�ߏ�C�{�Ï~�#�ü'����J~r�$����c�CF]�і��7��V�e��vU�F_�P��J�⌝�ʟ�݄m�TMNu�g�k�E�Ɓj^,}�9��L>�z�<H� ���FZ����7�).&c	�X�WyAS]�#XQ"Ucb�
y�y����C��Ct���#�+.�;)�c�>����[�o�_�}*Y�R�o���']F���X�ԓRP� ��^��͏J�¼s�k&�jod �����_�����Ð�}��`��<PO~+䞌�����1�כ�(���?.���Qyc��^ײ�6�^:9�܅b�@�(�z�[�j. �[�����e kLx`�f���N-uo(k/5nbK-�$�G�=��A�K��N�Q��{:�f�Ų�EQߓ�>
j½p�[XB��Z�@-�gX���u����MI���/�B��g����D�@��(} �]�V��9
�3���[���;��1���p4t�J6�E��E#��5��(es"d��>q�_#��j_�̜a�R���w�{T�W�͇?�a3�t}8jd���Y]-;���%���]u��M���p��W�(� ��|��A�í�x}(��hpȂm������0�({�Ϛ*�r�?�V�T/2S�FEp(D�b��𚸈��=^�Π��E��<(zAh�e�6F)�d|�����I����ڱ�A�����D�_�GJʟ��$eP��@%>(�8I��WD��͵���ͱO��fVO��V�Ŗ�R�fd�o�3�<7]SY����~�%�Y#�Zy`<��m��fc�^��k�u� MhgFf��yK��rke�+�Z��/^�r�/p��`<��ۥp�&D�%$&?�#�`��R@^���5�e�*l#��lb���>�*�U�Vc��-�֥ב��B�d��R<\JQ������^�F~�����Pl&/y##0�P��țsF�)l%Ũb*?~�@d���K�Y�v���&��l��ª����Q�@�t�t�b��+Ua������Gख़��gˀVV��f4��6���暊��z���sm��3����tq��W����V�~������R����uq6?��=��?�IG�&-����($��m6)E'%���>�z�>�.Z1�k��&G&�X�:�֑Gi
��@��>���}�/�]�\�ue1s��7�Z>���H����
e"�N�FU���0$����jH�Q��������1L��������<\�7m���I+��c�!/Y��pH�o���?��&a;o4H�3��a~�9�;ƒ�����FyzJ��#-*�Qa��s�O2q�~��W�IǺ�z/r~c�(H�,�}�))�)��G!yإ�<gx+�_�c�X0��؄��,�~eD��M�䔬���I�s\�dI�O�gAn��Ip>'�A�)�t=��gk������,�f��ZȔpTX��%�s���t�:�9'�!#�EC��z�#�����M�K?#�~�;JF�2589�]���,5lJY���Y�w���04�.�T��0����tTlQiz�uBz���jg�j���9���t�VR�Q��ku��ʴW���8�}�Qc}�V�����z)g%"�KO�UB���C�DV"x��+7����?
DI-����1��krj�q�b3-R��z�rC��5cA=K�ԑ͔��x:&ŏ9V�[H$��PD
1�D6��;j(�筧�{�~GAWh��=��A#��b]K���Q��(�;�<�&���`S�V�J�S�HcEH1�-���܄�Ac��W3=�~kԱ��fe�Q{���к�J3�߬·R�j8�a��ڪZ�IȔ��:-'O-B�db�zG�k�'��/�������ڷ��5����J $q$pa3��w��h��0)�=��::Owg���j�����5l�^i������2���#-*����^�h�q_�&���r�0���=e�g�CǪ�i���PЊ�9��E��YH�63^�o�;
����N��!;ϸpu���?d�,�t)�Q����@H�{�+]'��3؊95��0VA&Ǖ�sOZxձ/�0�E�;�.�nʍCc
�:�s�OǤ�u4�Oc��i���a�&�c��]w5*VU�z��Q�d78M�=Q�����h&��w���o�a��e��
ӣo�(�&�b�<� դUa����)�YY8R�,��$��ީ�gx,�����'/O�s&�
�
!�R&��QQ�����ߔ���(�z����^�+��<�Ƃ��p��<U�1�h|)�%e��������RE�'#�X��?�C���?olճ�uZ���e�]L���	՟�Z�9�:�����PP�'�Y{�4��	a�Y�������?�䨄>Jm�:ʝ��m7?���OJ��P�E���_V�x�]`�KC(�j۷y �}Κ+� �u)b �� �_~y>0&�:�.�&.�L���g6Pe�kA�v���,]���j�l����W������=TL�
�M�ܟJ�'�T�7�wW3"��b�0c�q�x� Y�Eԙ�c�#)�E~"D	LY���9yT�Dqr���sնx�׻���TG)�V��/��\�Ej�:�K.&x՛�!5M<G
�)�$���+�cW��y�ᤓV�=��==�J�7�m��Px�Ǭ����z�Ø�[XX�ɴW����]mC��3�8I����n����M�q5N3�==i,��U�BϬ��Y0���B~<�I�l 3�T ��&���Am1L\���Kp�f	[m_1��!��������O����b�^� �$��$/�Rca*����(�K�$����Q���E�(�F���R�0�S߂r�a(D! ~ON��2d���z�������﫝sJ�Y��XT���t����W�e1���{x�P��T���q���q$I��!r%[�jIX�d���z�<��p��ׇ+���NW7׫�<i���6��M���I$��N%��o�J]�d
��|����c��@�%�l�ޡo0~?��B�pË��v����D�&�?� Y%*�A��'� ��K���	ca���<|t��欣����u��ӻ�
oy�xkE@�[T� �(j��7����t|��b"EJU�A��X���D�U9	��(��Έ3�3�󂹧0k��TU,�w�qǍ���ʯ+4+��T��74&tnԃ��cn��؇�FOPV�+����ܳ�	'�8!�KI�˥Z��;�d|��q� �6�<�0�<��ʧV�cc[e(�ZCӗ��l	��>��/�ma��w�yG���_��}40�
;����V���?�~'R'7����&�,f�;�!�� 4lrtt�A�i�X"�e�w�.U�
��f�2�����lU�����
1�z
��(>�������M��SY�:&�z�F��>Wa+�����1I�,��_���S&�x!�B�SS�õ������4��&�����3��R��������[��ݏ?.|>��`���o��d�bU��v�iv�4����(s�'�|bڏ ����3���w�֬[�ſ|��ê'�O{�3�ҥ�����-^�]���Ӱnh��e�Z�%cc[�|�֝^�����љ��
+W=���DK�?t�l�bQG�7�p����Uk�QO?6��*�R����N-�<
Y�~Mz�bXF`�{sT���#耱EO�J�AU����G;,|�<����ĳ��8��"R��{x��d�VP�����E���d��ZBQk��W��ZBaފU�x�V�.��'�=m��&�E�|\��Y�F��ys�KKR/�m�������4W��|������}O���Ҽ	����V\��`Q�oi�R����/�{��a]T��w���9,�M}����~���p֙���S�@����([�ʴW��	@1���Ι3;U{�o��M��H�Kw�����?�)~��.�����}���?��!y��7c���z�^hȋO�y6YXF>��cͶ���#4�X4X��,⛅��
p�F�E*O�;ؤ�*\�7��d�Bl���a��yy��M+�UQ�D���J�
�H����"b!-g̞�{�y�Ɵ �����֬��p�C�5��r�~<�Z>^}������o��C�f_��O��p��[N�s�?�lI����
룞Y����_�bx�E�	wYl��#;2<�Уa<-�g���	tW��K���m
s�v�[n�U8���򽉟�5k��;	����as���zVX�nc�����z4�<� m!�x�	<4yx�^`�#{�'�MdYy���������O����C 5Ƚ2���h�d����^���tN�!:��]�"_Q1Vު�ڑ�$�����mC�WJ�U�L3�7�"2�\|ިH���0��[woC�	��d[9~�ܥ�{�dk���И���?�"�EO��^t���1�c98�F�0�U�m֪᷿�9��	a���>4d���ӈ���V�z<>�V>��z�r곭Q�A~�ӛ��F��Z�.ȴW�I#��RͲ�W���3<�أ)�H�ue-�Y��G��ąN�E �o����`g�y���TSx�'���/�5�җ�4��_�e���'ێ�j)�V�r�-,N��aq��M=�d[�SY|�{�e��D��?��Qdx����˛$L���ӱN� y���i�B����~���r�O<�8��
�%��@�+W��{�p��ˣ�9/.��3�� J�[�TaRl�J��<��,���.��#�?��p+���W���PO�B�ء,�����!+��������>��+Z!�ërχ|'�/I,P
,x~G�׿��f	(^���b���M�����+c���V8g\e�QԬF��9��'ק��L�թ��D�PR
��o�C���y
)��~����/.J��0�"O�WI+<Hn���%��+����}���Q�j�ĸ�GT��
�R�3�W:�EtpB�8�fu�����A�E���<�#�^����jQV�j�u��7����՟X�]�ܙ%]C�����qM�:�8�,wA=>a���ĘZ���7B�8U*�jB�4�!w+�˒Ŝ#�gC6�ERS=��E
��'baf,���~�|�m��62
�Qb#�0��&Y���IǦ� ���檼`<\B?��Q���+�'�=x-�a����\\l���e���`^w�Q���OL�uk���W��ು�ƥ����[ݳ���`�YJ%�!�^*u�M*UR^n"�{!atS�^���O��2�L�>�{���y��U�F�8�BGE�f�E���L�\�ĥ3�K^���O~Ұ� '�˼=e�A߶�GDʟP�^O���Cё����~fFA��B񵒱�C@�`
���G�&��	'�`s[ʜE�ӷ�������T�������ƅ�V6�r�_�V`��j�~{��.:�3�#
�&���L�z&}�tRp�kf�ww͊�¡��Fk}m�Y��h�f�QBgX�;�Ǯ�W���?�'}�Ї>d�>&(�?x j�۫ց�(�y*%�&+b4T!�K�[U�;j�E�����F��-*��)  �G90U$���J�W�J�z��b�Ó��]:v��!� ����Kx�0F�(:'e����9�ȧ���k��5���:u�9���u����-�bŊlA������UO�L3���	�j��O��]ʉ�3���{Pxr�C��G�aH��*�P����[������ ���Zgq�f�q��)��(8٧>��N)@�>	5��2��l'%(�O�xK��
�R[;�0QhB2�^�>�-��4��c,����\�\�o��2�h�񊮗�E4J���Q�V�}��P��u��4�p��>���'<��á .��]�E	�gO���ݢ�K�,��E��v0b^H��<M9"�T�_ٴW����#��}�s^�={��5�+,�.�~���~���Ҙyq�8���1ǝ:����V�V���
_��YU	"ڽa񫠊���<jH��2A�Of�_��2�t�bX�8����w�(�;��d�c�|��4变r���ɂ��fAP������@�I�&���������������}����k3 i;��cC�^{Z���ݖ��_���0ؿٸ�6m���ts�qǞ�v�3��p��	�@J��3*�g.�O�2��:+�B��������0{ޢ��!G�E��m�;V\n�.w5���h�@�I%7���d ��ӟ��n�����  ~� Ą(E�KJ����SF䕨���b�0����D������־�4�CV�����lq��
������A�|�q��L���D�w���	>=���¼{e��KϷ@�v���s��>Av��n
#z�~���1��%���·{ "��>!���Q�0>��������]w�i�Ϳ��?��N�,�T�` 1�1��$�İ/`�%M���G��M�
!�k�C�3�f|݊���wb��Sqt�d��zvO�O�����X��w��k�i�j�A%��aNT��.�?�x��E�=w���:��|�!)d��6n�W�ϕ�_c��]��{+3��O����K�f4��=[��Z3����h�����E�ȨU5��j�0�:���M�!\pAx��^��o�&\q��k_��YLLmW1Q�&k�S�>b�����K�"��k&n9^xb�hdbiۂ��կ!��j���I�ce��NQ��s£)�*�@�d#��+�b��c���$�}G�yOD��"+��'���WwM�P�B��E�+��B�B/�h��_�<�����@B8��������E�r�,
R�x�į/�����;�1�c����)��H�D�9�1����s���crO�f��o��`*����d�׊sa?P��M����4��/_ȋQ�󊗽܎o�Ż�9s���?$<s�)mC��>�9�P� І�%���)4�zjB)#�O�z֩,J�:_է�7��$(�!_@�]Y)bGT�NJ�6��`�Il����@r���>` ��\��p�r����0Y�-�˕U�;߃�.J��	Cų��H������{r�RZ:�S�B�Hd=QX��/R�οނQ�.�G�����ENVe=���}�zh��q0V�@*���+�}��Z�@,[�0�}�7�*c���£�������LfOx�P|��zECq�T�KIm�k�����~��_<�@;g#|G�~�Be��wA{H���CW�f�q.ox��E�C,<���/�\�1(P� ��K�~��~z8ꨣ�;Jx~)^3���/䞆�Ȍ%v�����WX��z�M7�
#i<ł��Z!��TYV�D����o?+�Fi��]v�e�\�w���h'E�+\�5�Ӕ2�I�q�9�+_��m˔t�:�!0�Aqބ��;����;L���t0�\�Rǣ�g�{˓�c����(���̹�]����X���z0Cmϓ�),e�C2��T u���gE��!U\ �u(�(�;�qSj-����3�Q��\s���/Xؾ�	�
�"�f������?�+Xy8@�Qp֭���	�O���Y �sl?ߕ{�x�o����g���O�$�'bM�}��,,X�Z��6�	p��싱��x���x򋱮�t��w,:��X���g�5C�Z��`�q=�y��F��Ɍ�zZ�Dq�
kEn�o�"�M��h���{��)��b|>
�N�@�L�`Q��m-��@�M���w�-&���x�O~�܂`���/�{�7V>��$

YҜ��d�� N��eeyŞW �}Ja).�܃����X����+9=�2Tx̋�ڢR��)T��o��d�_�t>~�-��Ň�t>�影Qצ�IP¬�Q��΢ �C]W�	{0�x-CB�E�Oޯ���<y}�7�a#o��Ʊ�m��x��[����2�ѥ������m�$�6ʱ��x ��?����{��^{�:�	�1�(��A�����9�ЖI����3~�G��c�'���C�EI=]\YA
mx������c4W	J���X�X*��b�a��O֤� S[;3�G�_)|3�'��%��%7ٷ{�y��XM����x��5X��GǨ��rqY[���4pM��G�z���U�P�6R�XO�c��ݓ+(�O��ׄ�qY�+�~�H<��,:)1�g���|2��̞~z,eQ�#��Z�-�~z����w��[�K
VcH��C�}���3�SCH��@ʠ�exCL9,>c�1t�����Ka�H}��G�t���9/�/0w��_��WٱC�v����X5�}N�/�X�bDe[\C�O��P�)%��6�><���ذO�q���|#����nAt�"�|q�@#%��.��P��J�MF�Y�?ɋ�d�MB���)��OhY%rk-ќQ:�[ ��z�%�BԾ��P-Z]�da!����?�SM���J����$X9f�l�� ���D0� ��x+�uU��{����Qܗ����a����l�+FΟI�dS�h��'Q�,��(/ΗEoO�J�EPJSR/���ל}���kxl��d趾��ay�׍k�}��5��uQ�����cD6�[J����!$��'�M
�Ѥh�țf�a5��߶��·	������K1yY�7�ٟ���;�7\3§�w>������w�Q��uև�Y�Q�Ωt�s�y7{�\�� �cp6�z��a�&��\`o�!B�ԋ��X�B<�#�G��� D���`>~�d�,���QP�E
PP7<�I>a+/AJD������}�Rg�qFn��!��J�Q���cb`��!�K����-������^JL��(Y�LL��e>���d��Zם�1�u�@��mOׁk&��~�m���|�3��/6����d
�Ca��C�0Iz^{@?�|���X
�#�|e�)<H�k�H8��
s� ���J����'��SO=�ƙ��
E�K��s���k���4�4�=�*���xd�(SZ�8O�����d�)��v�NT��%ijOpj��a�>8G��]�앰ւ�ךk���n@縵R��8�������U6�����2R�>��x���b� �()[M\�A9�*B2%KE�X�P���ؒU?9�ө���R*��� U3���ۿ5�Id�*�^�W���T��hC	̕���Q����(��4[�t<��|�+��ҹj��9�""h2E��#�J�^0J��9�z�ߏMY��������gD^'���'>a'��v�(k�G��vAa�X\r�%f�{�[�iy��7���"��BCR��X�}D<�Ya%b�,:��\�����{!EM��d29��H$�-��_�a'?������Y����Lsр&~��镧���y<dybrJ��5p������Ʊ�� ���#���N����{�]w�n�_ F�m�]n�$��R��`��*(~Vᕼ�}�3dぞ�J�+�Ȃ�� ��N*�=�n���9:�f��q~��"�?�S�I���V:V-��/�5�����%��-�j^���,s�÷��"� ��R�4%�j[v�裏��|��W�DM�g'�t���p�KɃ� D �������*�$i+�F2�y%wQt,v����{����o�KȊW�/��bJ� ϕx4��%����Dj#�6��^"�<���#EĘ�e�����'j��v)��\�;�5�\����CM�Da�Md��Z݊댧���
eP��"IG|]�p��y�"l�U)�c[�7ҙ�������X�BQ���R	b[�����A
�)�%�4��fA:6���Ci�UO��	��|�BB�7�Rj�����
�u�%n694h}�M�6�+��F������*�qP�O�KK�3�U-�_�1S�L��>mIe[c�8v�R%����ڗ{�g(
�~*[A�YӢJy���C@��e��Q6�3l,��k��������ߓ��WS��Nŏ$�����Ҵ7�(V-1H�C��U�XWL\�4)���~�����b�m����ZX�@�����(�w��?�m�Qm��(Y�L���,��s�U�3�����a@���E��1���Çu�:>�x�0�_,����\xα���y����D=T�T�i���{�_� T�3������^n�{_4�s�Ө}���Ry0�<N;�ܪ�ّE���J㷼�-�}�z�8�[��m�6Q�{"�` ����+_�J��!�O|߃�(���/�+����R����B-�����q��m`xlM/�F�P�^��TV�ȴW��=�o�!g�D�z�*��!FK�"b����CDV��T2�Α�,�?������\�h<��x-cS[ƖV8{Z:�H�׼�5�ȧ��<�*h՗ZL�(�������s��/��3Qt��G�ÃT�f�*�Y��yHo#)r yU������/	Q��2�?@'�����d�Ax�5��0�ô�s	���	5�:���B{��G!(�6؟&ߨ������6�,��a���>=����d�����o_�p͵�U�O�tWg�q������MZr ����+?&D�i��&؃���[[W�R����B��b4<h|M~������X2�Ǌ_(���
K�"����`�\��j[������(�ָ}Cx�����k�r�=N��y b�_08Ny�~�C'|~�G��A�!Z T9��=��XX�,>$�	E��R����G���������Sjܔ��Tf��/%;�寄����!zx%!b��Jx�b?ȥT��e���-�&�`z��9���"���B�!o����G����.E1���6a�f���bbX���)���R��<Q��W%F��4O��b&���������o��
ay"E_��{,���C*�!���������X����u�[��Vر�xE�%�N+�B�o�<�?F`؉E�@�T��^
����ʁ+�䘚ë+������9dWPȂb����rDC��[c�f��I��}c�q�>o��V;z��H�n7�0��m$�ے���3x. H��o�h�IE�+���}�E�����ٶZ�"���V�%�g�D���E��_�%j\� 
���k^͇<���rQ����+�s�8�����M\vV�ǟ���ʿh��l7Ӈh'[!,!^snX_|���'�{<N�X���˲?��g���|vu�\G�F�o�zƭSA�=�xA6Fs��E���7��DSma�;�!h&r�Ց�S;p}��s�?�g[R�u��1(G�X��ͮ� �,�,�(Y�� �4��<+�((*�����18 ��,�Z %�C~�Lh��&d�3���2ɇ)?��T���(�ڷ���ۙ%���TM{��lugV���n�s)��9_Q�X'
Z�Lաk�I
���iʚm͝=ǬtQ8�j:=�����r�-��ũ�dR<ZU���X�g�u�uR"�� ~x��!�Z�#+�,Ă*ب�rK�E`��/Xo�Ḋ���U�3ް�?��O�7�����_��_�؅�����YX�4Ua|���4�-�U^$h1�Gq4)���2��1I:�!��7F�ƫX8U�"�-Q��z�m≰�����_)猻;��k�TJ����������Q|��^���M_��}�K�o\V\]�$s�`�z��>���d��
b)
��@Lo��f��O,�F�����!V��a7�/y[=g�IQ�y=�>��R�x��IֻN��#Dm�X��(.:tѪ%���7�$���XM�W�1n̂��@�?1��lC�Xǀ�[�2�+'����u��	H&���DH�?IGwG��ŴW�q�k��������I%����'��-Z�>���dՖ��N%ٔ�U��1}�6D��Ќ�5�W��U�Țc1�dl$�0<��9�Q��W�V�~݄�����L�o$j��ppO�N�?��8��҇�9�I��C��#���F�TM�Xt�z̿��=�� lKy.O�k�&C�J�<Ť�3��.�b�?�fo�K�B.�X�r�5i4@}`O���C���)���7�֢��M����ĵ���\CV�g�(�3AU��X�R^����D�阽���,E˾���S�Һb2k��ux�8�h���W�D�"P�9�43 CUOy �k�Lݷ<�ƷBA2<|����YO���VD��+#�-wf�T��==s���ٴW��Ty�[�^	*�3�E3$#�gE.M�9����D�)�llk�%!�����xeQ��E֥�s��e�Y~!Cl���6��˛%�&�/
�
����+<!k��J����\C*TI(*	�1#��S��s~?���י�&	UOR���:��"f�b=�>�\�:O�_a��G��O+���U;Ey�y&zD����n ���$��Z��K#�?U��E4n��"���_{?G4�$;��/gƛBV�����{.YR� �ښod�����7͟?��M�Ԓdf��+��H�Q���׾6\t�E�$D��r~��sP <�LEbp���z��$�'��T����b"���7��h9u@Sӟ��!�g�#��8F���Y��9%�E�,�&�4�t}�U�:MT��<:mp�����\�׽�u6>�؅n^���ã�?6�8i�։<o�5����ق�n�=������O��{�d�ƍ��w�&�T���D�&%���Lpoa1�9a���Ț���@�(!rI��	���g��_�z����R)ԉTVń�Be`�9,y.$79~�!�bƱ�:Y!���3Q�L�+��W��ն/q�����h� ����7j���˾�e�m�ehK#Q"]p�Y�O~��+��v�+���-��Z�7^�C�"k˶��1`���y�ؼ����b��C��v)U�i17�p���k� CNm�JHM,A'�'�^��c�'�������
˱ `q�|W��^��(�a����J"��K/5���������}�5�� ��7����>6�����!�EcY9�ٳf�{��'�-Ӟ�����O��v�i���\��5ض�'f[FD�F5�'!t��=R�R������ʿ��  �IDATK|<_}x��Ǫ�E����C$F[BO�ࡒ%EZc�&�΢0�^Z�|�J�m�d	��ZQ��9��0|��9F��.��2k���9v ���+̪�C߄�[{N�.�gK�-���u�p��ϸ�W}��o���GN?���]u��/]�p��(+� �k˶��v�!t���A��4)N�EL��_Oi��P%�s�,F*�����{,dB�����o�=��_,�B�������*����.�U���eL	j) <�n\S��e�b�E��G޺�0��x[K���CG<�w���������W+N:��xa�V����.�BJ8*$E]J�����x$�^���#Z8>
�(tCD1�r����%�&%E̽M%��P�6���
�����VHj,%:Q��J|q�GSi��?���jKt���el�H7�`�{/[��?��?�g����~��߽�_?;��T�����˷'[�dbЩ��j�	��LLe�'��)&�z�h�Dr��5�����)�9L�xxa���'^W��ؿ�f��F�Χ�5�����ب�=��S�s�i��q�����ZX5�5DiKs��F�E���U�|�W�n�(�s^�������>��p��܍��L�3�҇z���r���1�})
D� ̻�cҲ�FB#F���g�T�����"��p���#<�J�[����2�$�
u���CY�r�J�������dm�߱@;}���>8g!l��6������p.)�^�~_�s@	�j����}{�"�Aq�~#�c��)�(rA0��]�a}8��s�Yg��~[.��,�_����}g	ܡ�P��W�@��ZĔ+R�]�FW�.uƶƱ�PZ���:-ORM��S�ҟ�\������ ����贿��~�zvϬ[�;�[�v�(���E�\x�_������y!����3n���������Y)�XNr�Q�ziԓC���'V>�+ioU�m�(�,w~���z֞��K!�G0V�/v��C\K���?��k���J��x�a��^���:�!X���ndyRؾ�I!�祰�/L���J��gG������Gы�Mֺ�N�C��Їrg%�=lјѽd~�}������^DcQ�V
�=�P�M��>����<~�,�>G��Fk�#�2e�{ Bu��2��5����.�����6� 9�S���{^o�y�Oc��^��d��j5�h��"��ui��a`���:�+�f��"~�_�x /�1���+W�H1�>Q�)7�S�� �}ݚ����Ś���G�Ņ�,��x��\��r�0-
Z@����/�rjF�_�=�_�I��2�����A�؁x-z_:N]#]��H����s?���=#&"h,�џA���C��gh|	��חmiAW1"�)�HV�Կރ��G��M7ݔ�85o���}��;�h�^1��8���/~�w>��4�݌R�тz��o~�7�x�aq@h�0=��Y1�~D�O�q���R��)��&�,:Y>�z�]�c*���v�R�2(�B2J&2�e]�-��yJB��Q�C�аV=V˵�-�~~�P���Y�=�s`�{�+^a�y0�:�΅B4�g�������0��̈́��,jfy��q�������*�H�PD4��Aޙ@��}���c�,7VaZh�D�x�Ɍ�Y���&|}�T塘�5���C��3�<���og��G.���?��ˢ����'Ƈo�T�鞙����Wq�vu��1֎�&U��\<�rɬ�v��L�<=l��ΏG��~���&�b�b5�����6����{�"�_�I�&��5���-=����
���h��G<��o�鷃�Z������J$��B4�Z0u���4v���Tϓ.BZ=��b�ڎ?�/�k�,�d���l�"_F�����4ߢ�A{�0٩*Zp�O�Hظ�{|����[��S�q���?�㣟�������%Qyv�϶�?O� �#7��S��DO���\T�|�Ᏺ��p��h��Q���G��w�����xp��U�+�h�vw��C��Z-�,�Ks�RZ�aÆ���^��D��v*�k%���TW0^��r�|}��DI���¥~(~y���=%c=ݶ����B.�7n���v�/Nd%�Y���Z.��̍����0v ��xF_��+dO��Yq�Iy�B4iq��i�>�����@Ź,c�'�=/�S]��ո@��q���.�<��ȌS���_���~������V�`�EG�B��ʯ��OZjB�
�sd��z���'�����)��p���|�q�-#):�����̙��W��e�~����c��c)'=IG)�UX����k�w*)���&�Ox*<!�89!!W`�$�O')�<�W�zo�����!�c�9��9�~�Y�
�(ɫs�sy ���/��/_~�G?��w�m���<^��ZT��4 ���X��.��ҷ$õ?�;{�"����:�dF�g-zr�XK}�L�^cYqx�'�����1���Nr�_����h�X1�1�O,�����/|w��[��T���_�����߿��7\s��M�o�T��RXr�YU��M$}֊����2�a�714�O<?�(������q=��������o�г���Uc���]PH�k��{�`m�+$,W�IAR�bŊ�ɷ��,h%=�7�=ďC�p������V�C笐�^�|��7��y�I'���&��骫�z�%�\�!n�q���1d^h�����},_�(�䓻S�D����g��[^��x����/�QP`-�B�y0����P�ђ|���{sl�og��G����7��w�m��6�n:;��]
�zqmo����+�O) ?�䎓��i�mb,��b�԰�jõQ
�Oબ�q��5�dg�GY�x�_�����G�R��0~/#������>��Ǉzd�J���RH�ڄ��zƆ���?��?�Qu�x��Op���;��7\{������x^�c���șI�
e�=���O����ւVTƾ���-��Iw�������]-J��9}�y{���j���6Z��L�D�B���*����y�����[�����~�����-oy�O��M��^T��R����
�Qp�V���sl�뮻.�p��H{����I��W��"���o�#��څ�כ����x�O4���81���>�+���L��^#����Tq��vi��9�3�_y啗���kg<����4+U��\A�+��зU<�����pǈ�{�ޒ�I�W3Δ��h�f�;�!��� FyGq����֊�W\������n˾g��G�K�ȥ��M���OƋ��Ύ��!�Rф:T���PK�\&Kd�kr0@�!x���p�
	��Ysf��j��;n��N�O�&Չ�+tuu�[�[���w�p�	<�y��{��8P�[a�}��YR��r���a���	����7��E[s,�{���/������*q��׻��X�2�a�l�h;��*�v����z��oG����9.���줮'��kL����d��'-��������u�kf �)m�ɛ_��W\q�;���/���G~�O��d~��#'d)7��<���x|AS�2�
u�}&.5��"��Xg���)/�XY'��/���:�c�)~N��؞����}r\q�f��tW�^+�-Z��YO|wQj�$�?��u�\s�����q^����W�σ�+���(K��m(�������#$R����d��z��>
�f������M�q�^�]y�Ag���l+'�w�����y�{����\saT!�tw/����Cx�f�{{����ng�q�s�����y��Y�U1�r#�6�Y4;�fʩ�ҁ%�v�����+_�J�c���8;�.��{�0fY��9�����<�Fֲ���!ت��n�������:{������+�,����#������^�|���H!-e$��x�\&���*e�|R�I����h�<�`���8a�G��w����}n��n+�:��������ݯy�k�sϽ��q(ύ7�8��;Z�'���|��P��^\����M����m�������ۗ/����u�Y���ٽ��.�&�&s��=��me��]<��O?�l�n���mrmN?��M�������O��O�|����&"i�p���P:R���h㦈������1�&������=��1������ӎ���ۿ���+���}�����?+ޭ�{�����7���#������{��7g�x�:';��	�T��	���|�é%�QU�B�H�5I��3�C#�+_��׿+Z�+C��z��Z�kD����+��s)�����a!FY�8�c��ړa,�����>���;����x��ZI��"���7�a��o=����-�&W4�8&<�x�6Ɨ���g�]��O������{����	�w[�� o{���>���~��{�%��y�Q����dxy\v���0]���WI$CV~R*���L.8����YSa��JI�aҷysR��`F��,,g�rV
S.�=���R*ل��;R�YRuk�4�`pB��RP��;E%b�����y�m���@���x�?�;g�G�F�#��wߓO<��/�.]J�w��Y�f͉(�6'������q(��bի�#Wz���z��Fp�Xyka��%�F����x��h�sSk���^o�F�go����9ȧz�Wuu^�ˮq��R�G�X;���@�}��J�8G������m'ʽUʕ�;*b���Qf����8�x惵�����rg�(���R�RI�zŗꎇ�}����'�\J[ܛ�{T����j_<��{�������C:�8����7��(m�������W]uUwTB��гf͚Yq0΍�DԡS8�y\��%j%dcJ�n��f+��w������7�3N�2Ǥ��5Ǥ��/����&�4��1��uR��'������~v,���qL|���K�������x�~W�Egէ>���ƒ�x≏���?�hT������R��n^�#�e�m��3>*<w�7�d��g�W��H���Low<^����.���,����w	r]�d�Prz�K��^Jo���&��4����@��@�����uB3�;�Z�T��{���;z�I��ܶ�1�W�XfPƱ�~�u����gOs�1�V.��~z�;����y��ٳg/�ے���.u-;^�A5~n��{:���������k6��㸩e�|>_�h��yvM�l��`���K�=*�����54��M�D�%��&��9r<�cw .��K�,�׭wٲek�9���7�%m�?9�l˶�
m��r�i�Q�{O�d�&�(o*������k��Z�%�z׻n�nm٩����ҖqH�M�J�������[�Җ��@i+����-m���V�miK[�2����Җ��eJ[���-mi����oK[�Җ(m�ߖ���-3P�ʿ-miK[f����^��2�R    IEND�B`�PK   �eX��=�)  �     jsons/user_defined.json���n�8�_�еipx�����u�m� n�
��$*֖T6�{)�*�-Q����3�<�c����kt�=�Y^�4�������<s���~h\}{:�Y�]���ꆒ�F7����Vߕ��|5���Iv3�ԌϨ̔#�Aq��H�Z!�H	'�^��Ue��v}��yֻj�N?�l���Ϋ�8�ˌo���'
CJI�T�%b*�(&R �!�@BJ0L���<�'eq|(K3��(�,A,��d(#�NC�����N�鏥Y���5?����ks�ʋE����SPt�Y�T[�8-�f7�,�3�r�|��21�"�(q����tfU�"]�un�F�P6y��o�+��$bL��`�iOț��侬����ۚ��X�p��^����M?S�� � �pO���\ � V}��'��ӏ�X�}`?b�ҏ|��U?t�K�V@� �&�V�t��`RpF���";*��+iG8�����rfG8�x'b�H����2n�u���i�5��ik��5�g>p:��M���6���+���&�����th틾�릟� Cc_ �%�~dh���q��=�����w��
��� �K�#���������EC;_ �E�^�����%�"J�^~A�.���"@\V�/��^�����5��C����_B�=������:v��g�:��h�.C{����pڻz�n� ���k�c.C{WN�v����ỿ�������؍x�k�}�7���u���~
�[�hu���붭USy2Z�)�_����ھ�p�ġ)�*����!J!	Q�R��PRE�ցg�A�Ri,�Q0ZB����:�>����pr��u�HJ�[��a�
	�P0�e�j�°�-��N�/M��W�"dV�__^o�w��i���Ϩ߲�����t�a����8�x�ӹ����L�!����ᦶ]�ou�D���O�L�=E�}�𹘖����:o�x�����Gw�ΰ_����.SI�պ~	�T���]�؛�}�H-�����)F$#�yG�:�a��wsm���PK
   �eX	r+�  �Q                   cirkitFile.jsonPK
    eXǐ]zd� K� /             �  images/2a01d32d-a809-4abe-b296-5e1ff191d201.pngPK
   �eX����H   C   /             �� images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   �eX��) oj /             *� images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
    eX@��)  /             ��
 images/fdf90566-ce4c-4b91-9798-b6c065370fb3.pngPK
   �eX��=�)  �               
� jsons/user_defined.jsonPK      �  h�   